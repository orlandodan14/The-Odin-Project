--- !ruby/object:Game
misses:
- e
guess: e
progress:
- "-"
- a
- "-"
- "-"
- "-"
- "-"
- "-"
- a
guessed_letters:
- a
dictionary:
- |
  Aachen
- |
  Aalborg
- |
  aardvark
- |
  Aarhus
- |
  Aaron
- |
  abaci
- |
  aback
- |
  abacus
- |
  Abadan
- |
  abaft
- |
  abalone
- |
  abandon
- |
  abandoned
- |
  abandonedly
- |
  abandonment
- |
  abase
- |
  abasement
- |
  abash
- |
  abashed
- |
  abashedly
- |
  abashment
- |
  abate
- |
  abatement
- |
  abattoir
- |
  abbacy
- |
  abbess
- |
  abbey
- |
  abbot
- |
  Abbott
- |
  abbreviate
- |
  abbreviated
- |
  abbreviation
- |
  abbreviator
- |
  Abdias
- |
  abdicate
- |
  abdication
- |
  abdicator
- |
  abdomen
- |
  abdominal
- |
  abdominally
- |
  abduct
- |
  abduction
- |
  abductor
- |
  abeam
- |
  abecedarian
- |
  Abelard
- |
  Abenaki
- |
  Aberdeen
- |
  Aberdonian
- |
  Abernathy
- |
  aberrance
- |
  aberrancy
- |
  aberrant
- |
  aberrantly
- |
  aberration
- |
  aberrational
- |
  abetment
- |
  abetter
- |
  abettor
- |
  abeyance
- |
  abeyant
- |
  abhor
- |
  abhorrence
- |
  abhorrent
- |
  abhorrently
- |
  abhorrer
- |
  abidance
- |
  abide
- |
  abider
- |
  abiding
- |
  abidingly
- |
  Abidjan
- |
  Abigail
- |
  Abilene
- |
  ability
- |
  abiotic
- |
  abject
- |
  abjection
- |
  abjectly
- |
  abjectness
- |
  abjuration
- |
  abjuratory
- |
  abjure
- |
  abjurer
- |
  Abkhazia
- |
  Abkhazian
- |
  ablate
- |
  ablation
- |
  ablative
- |
  ablaut
- |
  ablaze
- |
  ableism
- |
  ableist
- |
  abloom
- |
  ablution
- |
  ablutions
- |
  Abnaki
- |
  abnegate
- |
  abnegation
- |
  abnegator
- |
  Abner
- |
  abnormal
- |
  abnormality
- |
  abnormally
- |
  aboard
- |
  abode
- |
  abolish
- |
  abolisher
- |
  abolishment
- |
  abolition
- |
  abolitionism
- |
  Abolitionist
- |
  abolitionist
- |
  abominable
- |
  abominably
- |
  abominate
- |
  abomination
- |
  abominator
- |
  Aboriginal
- |
  aboriginal
- |
  aboriginally
- |
  Aborigine
- |
  aborigine
- |
  aborning
- |
  abort
- |
  abortion
- |
  abortionist
- |
  abortive
- |
  abortively
- |
  aboulia
- |
  abound
- |
  about
- |
  above
- |
  aboveboard
- |
  abracadabra
- |
  abrade
- |
  abrader
- |
  Abraham
- |
  abrasion
- |
  abrasive
- |
  abrasively
- |
  abrasiveness
- |
  abreast
- |
  abridge
- |
  abridgement
- |
  abridger
- |
  abridgment
- |
  abroad
- |
  abrogate
- |
  abrogation
- |
  abrogator
- |
  abrupt
- |
  abruption
- |
  abruptly
- |
  abruptness
- |
  Abruzzi
- |
  Absalom
- |
  abscess
- |
  abscessed
- |
  abscind
- |
  abscise
- |
  abscissa
- |
  abscissae
- |
  abscission
- |
  abscond
- |
  absconder
- |
  abseil
- |
  absence
- |
  absent
- |
  absentee
- |
  absenteeism
- |
  absently
- |
  absentminded
- |
  absinth
- |
  absinthe
- |
  absolute
- |
  absolutely
- |
  absoluteness
- |
  absolution
- |
  absolutism
- |
  absolutist
- |
  absolutistic
- |
  absolutize
- |
  absolvable
- |
  absolve
- |
  absolver
- |
  absorb
- |
  absorbable
- |
  absorbant
- |
  absorbed
- |
  absorbency
- |
  absorbent
- |
  absorber
- |
  absorbing
- |
  absorbingly
- |
  absorption
- |
  absorptive
- |
  absorptivity
- |
  absquatulate
- |
  abstain
- |
  abstainer
- |
  abstemious
- |
  abstemiously
- |
  abstention
- |
  abstinence
- |
  abstinent
- |
  abstinently
- |
  abstract
- |
  abstracted
- |
  abstractedly
- |
  abstracter
- |
  abstraction
- |
  abstractly
- |
  abstractness
- |
  abstruse
- |
  abstrusely
- |
  abstruseness
- |
  absurd
- |
  absurdism
- |
  absurdist
- |
  absurdity
- |
  absurdly
- |
  absurdness
- |
  Abuja
- |
  abulia
- |
  abulic
- |
  abundance
- |
  abundant
- |
  abundantly
- |
  abuse
- |
  abuser
- |
  abusive
- |
  abusively
- |
  abusiveness
- |
  abutment
- |
  abutter
- |
  abuzz
- |
  abysm
- |
  abysmal
- |
  abysmally
- |
  abyss
- |
  abyssal
- |
  Abyssinia
- |
  Abyssinian
- |
  acacia
- |
  academe
- |
  academia
- |
  academic
- |
  academically
- |
  academician
- |
  academicism
- |
  academics
- |
  academism
- |
  academy
- |
  Acadia
- |
  Acadian
- |
  acanthi
- |
  acanthus
- |
  Acapulco
- |
  accede
- |
  accedence
- |
  accelerandi
- |
  accelerando
- |
  accelerate
- |
  acceleration
- |
  accelerative
- |
  accelerator
- |
  accent
- |
  accented
- |
  accentual
- |
  accentuate
- |
  accentuation
- |
  accept
- |
  acceptable
- |
  acceptably
- |
  acceptance
- |
  acceptation
- |
  accepted
- |
  accepter
- |
  acceptor
- |
  access
- |
  accessary
- |
  accessible
- |
  accessibly
- |
  accession
- |
  accessional
- |
  accessory
- |
  accident
- |
  accidental
- |
  accidentally
- |
  accidently
- |
  accidie
- |
  accipiter
- |
  acclaim
- |
  acclaimed
- |
  acclaimer
- |
  acclamation
- |
  acclamatory
- |
  acclimate
- |
  acclimation
- |
  acclimatize
- |
  acclivitous
- |
  acclivity
- |
  accolade
- |
  accommodate
- |
  accompanist
- |
  accompany
- |
  accomplice
- |
  accomplish
- |
  accomplished
- |
  accomplisher
- |
  accord
- |
  accordance
- |
  accordant
- |
  according
- |
  accordingly
- |
  accordion
- |
  accordionist
- |
  accost
- |
  accouchement
- |
  account
- |
  accountable
- |
  accountably
- |
  accountancy
- |
  accountant
- |
  accounting
- |
  accounts
- |
  accouter
- |
  accouterment
- |
  accoutre
- |
  accoutrement
- |
  Accra
- |
  accredit
- |
  accredited
- |
  accrete
- |
  accretion
- |
  accretionary
- |
  accretive
- |
  accrual
- |
  accrue
- |
  acculturate
- |
  accumbent
- |
  accumulate
- |
  accumulation
- |
  accumulative
- |
  accumulator
- |
  accuracy
- |
  accurate
- |
  accurately
- |
  accurateness
- |
  accursed
- |
  accursedly
- |
  accursedness
- |
  accurst
- |
  accusation
- |
  accusative
- |
  accusatory
- |
  accuse
- |
  accused
- |
  accuser
- |
  accusingly
- |
  accustom
- |
  accustomed
- |
  acedia
- |
  acerb
- |
  acerbate
- |
  acerbic
- |
  acerbically
- |
  acerbity
- |
  acetanilide
- |
  acetate
- |
  acetic
- |
  acetone
- |
  acetonic
- |
  acetylene
- |
  Achaean
- |
  Achates
- |
  Achebe
- |
  achene
- |
  Achernar
- |
  Acheron
- |
  Acheson
- |
  achievable
- |
  achieve
- |
  achievement
- |
  achiever
- |
  Achilles
- |
  achiness
- |
  achromatic
- |
  achromatism
- |
  acidic
- |
  acidifier
- |
  acidify
- |
  acidity
- |
  acidly
- |
  acidness
- |
  acidosis
- |
  acidotic
- |
  acidulate
- |
  acidulous
- |
  aciduria
- |
  acknowledge
- |
  acned
- |
  acolyte
- |
  Aconcagua
- |
  aconite
- |
  acorn
- |
  acoustic
- |
  acoustical
- |
  acoustically
- |
  acoustician
- |
  acoustics
- |
  acquaint
- |
  acquaintance
- |
  acquainted
- |
  acquiesce
- |
  acquiescence
- |
  acquiescent
- |
  acquirable
- |
  acquire
- |
  acquired
- |
  acquirement
- |
  acquisition
- |
  acquisitive
- |
  acquit
- |
  acquittal
- |
  acquittance
- |
  acreage
- |
  acrid
- |
  acridity
- |
  acridly
- |
  acridness
- |
  acrimonious
- |
  acrimony
- |
  acrobat
- |
  acrobatic
- |
  acrobatics
- |
  acromegalic
- |
  acromegaly
- |
  acronym
- |
  acronymic
- |
  acronymous
- |
  acrophobia
- |
  acrophobic
- |
  Acropolis
- |
  acropolis
- |
  across
- |
  acrostic
- |
  acrylic
- |
  actin
- |
  acting
- |
  actinic
- |
  actinide
- |
  actinism
- |
  actinium
- |
  actinomycin
- |
  action
- |
  actionable
- |
  actionably
- |
  actionless
- |
  actions
- |
  Actium
- |
  activate
- |
  activation
- |
  activator
- |
  active
- |
  actively
- |
  activeness
- |
  activism
- |
  activist
- |
  activistic
- |
  activity
- |
  actor
- |
  actress
- |
  actual
- |
  actualities
- |
  actuality
- |
  actualize
- |
  actually
- |
  actuarial
- |
  actuarially
- |
  actuarily
- |
  actuary
- |
  actuate
- |
  actuation
- |
  actuator
- |
  acuity
- |
  acumen
- |
  acupressure
- |
  acupuncture
- |
  acute
- |
  acutely
- |
  acuteness
- |
  acyclic
- |
  acyclovir
- |
  adage
- |
  adagio
- |
  adamance
- |
  adamancy
- |
  adamant
- |
  adamantine
- |
  adamantly
- |
  Adams
- |
  Adana
- |
  adapt
- |
  adaptability
- |
  adaptable
- |
  adaptation
- |
  adaptational
- |
  adapter
- |
  adaptive
- |
  adaptiveness
- |
  adaptivity
- |
  adaptor
- |
  addable
- |
  Addams
- |
  added
- |
  addend
- |
  addenda
- |
  addendum
- |
  adder
- |
  addible
- |
  addict
- |
  addicted
- |
  addiction
- |
  addictive
- |
  Addison
- |
  Addisonian
- |
  addition
- |
  additional
- |
  additionally
- |
  additive
- |
  additivity
- |
  addle
- |
  address
- |
  addressable
- |
  addressee
- |
  adduce
- |
  adduceable
- |
  adducer
- |
  adducible
- |
  adductor
- |
  Adela
- |
  Adelaide
- |
  Adelbert
- |
  Adele
- |
  Adeline
- |
  Adenauer
- |
  adenine
- |
  adenoid
- |
  adenoidal
- |
  adenoids
- |
  adept
- |
  adeptly
- |
  adeptness
- |
  adequacy
- |
  adequate
- |
  adequately
- |
  adequateness
- |
  adhere
- |
  adherence
- |
  adherent
- |
  adhesion
- |
  adhesive
- |
  adhesively
- |
  adhesiveness
- |
  adiabatic
- |
  adieu
- |
  adieux
- |
  adios
- |
  adipose
- |
  adiposity
- |
  Adirondack
- |
  Adirondacks
- |
  adjacency
- |
  adjacent
- |
  adjacently
- |
  adjectival
- |
  adjectivally
- |
  adjective
- |
  adjoin
- |
  adjoining
- |
  adjourn
- |
  adjournment
- |
  adjudge
- |
  adjudgement
- |
  adjudgment
- |
  adjudicate
- |
  adjudication
- |
  adjudicative
- |
  adjudicator
- |
  adjudicatory
- |
  adjunct
- |
  adjunctive
- |
  adjuration
- |
  adjuratory
- |
  adjure
- |
  adjust
- |
  adjustable
- |
  adjuster
- |
  adjustment
- |
  adjustor
- |
  adjutancy
- |
  adjutant
- |
  adjuvant
- |
  Adler
- |
  Adlerian
- |
  adman
- |
  administer
- |
  administrant
- |
  administrate
- |
  admirability
- |
  admirable
- |
  admirably
- |
  Admiral
- |
  admiral
- |
  Admiralty
- |
  admiralty
- |
  admiration
- |
  admire
- |
  admirer
- |
  admiring
- |
  admiringly
- |
  admissible
- |
  admission
- |
  admissions
- |
  admissive
- |
  admit
- |
  admittance
- |
  admittedly
- |
  admix
- |
  admixture
- |
  admonish
- |
  admonisher
- |
  admonishment
- |
  admonition
- |
  admonitory
- |
  adobe
- |
  adolescence
- |
  adolescent
- |
  Adolph
- |
  Adonai
- |
  Adonis
- |
  adonis
- |
  adopt
- |
  adoptable
- |
  adopted
- |
  adoptee
- |
  adopter
- |
  adoption
- |
  adoptive
- |
  adoptively
- |
  adorable
- |
  adorableness
- |
  adorably
- |
  adoration
- |
  adore
- |
  adorer
- |
  adoring
- |
  adoringly
- |
  adorn
- |
  adorner
- |
  adornment
- |
  adrenal
- |
  Adrenalin
- |
  adrenalin
- |
  adrenaline
- |
  Adrian
- |
  Adriatic
- |
  Adrienne
- |
  adrift
- |
  adroit
- |
  adroitly
- |
  adroitness
- |
  adsorb
- |
  adsorbable
- |
  adsorbent
- |
  adsorption
- |
  adsorptive
- |
  adulate
- |
  adulation
- |
  adulator
- |
  adulatory
- |
  adult
- |
  adulterant
- |
  adulterate
- |
  adulteration
- |
  adulterator
- |
  adulterer
- |
  adulteress
- |
  adulterous
- |
  adultery
- |
  adulthood
- |
  adumbrate
- |
  adumbration
- |
  adumbrative
- |
  advance
- |
  advanced
- |
  advancement
- |
  advancer
- |
  advances
- |
  advantage
- |
  advantageous
- |
  advection
- |
  Advent
- |
  advent
- |
  Adventist
- |
  adventitious
- |
  adventure
- |
  adventurer
- |
  adventuress
- |
  adventurism
- |
  adventurist
- |
  adventurous
- |
  adverb
- |
  adverbial
- |
  adverbially
- |
  adversarial
- |
  adversary
- |
  adverse
- |
  adversely
- |
  adversity
- |
  advert
- |
  advertise
- |
  advertiser
- |
  advertising
- |
  advertize
- |
  advertorial
- |
  advice
- |
  advisability
- |
  advisable
- |
  advisably
- |
  advise
- |
  advised
- |
  advisedly
- |
  advisement
- |
  adviser
- |
  advisor
- |
  advisory
- |
  advocacy
- |
  advocate
- |
  advocation
- |
  advocator
- |
  Aegean
- |
  aegis
- |
  Aelfric
- |
  Aeneas
- |
  Aeolia
- |
  Aeolian
- |
  aeolian
- |
  Aeolis
- |
  Aeolus
- |
  aeonian
- |
  aerate
- |
  aeration
- |
  aerator
- |
  aerial
- |
  aerialist
- |
  aerially
- |
  aerie
- |
  aerobatics
- |
  aerobe
- |
  aerobic
- |
  aerobically
- |
  aerobics
- |
  aerodrome
- |
  aerodynamic
- |
  aerodynamics
- |
  aerometer
- |
  aeronaut
- |
  aeronautic
- |
  aeronautical
- |
  aeronautics
- |
  aeropause
- |
  aeroplane
- |
  aeroponics
- |
  aerosol
- |
  aerospace
- |
  Aeschylean
- |
  Aeschylus
- |
  Aesculapius
- |
  Aesop
- |
  Aesopian
- |
  Aesopic
- |
  aesthesia
- |
  aesthete
- |
  aesthetic
- |
  aesthetician
- |
  aestheticism
- |
  aesthetics
- |
  aestival
- |
  aestivate
- |
  aetiology
- |
  affability
- |
  affable
- |
  affably
- |
  affair
- |
  affairs
- |
  affect
- |
  affectation
- |
  affected
- |
  affectedly
- |
  affecting
- |
  affectingly
- |
  affection
- |
  affectionate
- |
  affective
- |
  affectively
- |
  affectless
- |
  afferent
- |
  affiance
- |
  affidavit
- |
  affiliate
- |
  affiliated
- |
  affiliation
- |
  affiliative
- |
  affinity
- |
  affirm
- |
  affirmable
- |
  affirmant
- |
  affirmation
- |
  affirmative
- |
  affirmer
- |
  affix
- |
  affixation
- |
  afflatus
- |
  afflict
- |
  affliction
- |
  afflictive
- |
  afflictively
- |
  affluence
- |
  affluent
- |
  affluently
- |
  afflux
- |
  afford
- |
  affordable
- |
  affordably
- |
  afforest
- |
  affray
- |
  affright
- |
  affront
- |
  affronted
- |
  Afghan
- |
  afghan
- |
  afghani
- |
  Afghanistan
- |
  aficionado
- |
  afield
- |
  afire
- |
  aflame
- |
  aflatoxin
- |
  afloat
- |
  aflutter
- |
  afoot
- |
  aforesaid
- |
  aforethought
- |
  afoul
- |
  afraid
- |
  afresh
- |
  Africa
- |
  African
- |
  Africana
- |
  Afrikaans
- |
  Afrikaner
- |
  Afrocentric
- |
  Afrocentrism
- |
  Afrocentrist
- |
  after
- |
  afterbirth
- |
  afterburner
- |
  aftercare
- |
  afterdeck
- |
  aftereffect
- |
  afterglow
- |
  afterimage
- |
  afterlife
- |
  aftermarket
- |
  aftermath
- |
  afternoon
- |
  afterschool
- |
  aftershave
- |
  aftershock
- |
  aftertaste
- |
  afterthought
- |
  afterward
- |
  afterwards
- |
  afterword
- |
  afterworld
- |
  again
- |
  against
- |
  Agamemnon
- |
  Agana
- |
  agape
- |
  Agassiz
- |
  agate
- |
  Agatha
- |
  agave
- |
  ageing
- |
  ageism
- |
  ageist
- |
  ageless
- |
  agelessly
- |
  agelessness
- |
  agency
- |
  agenda
- |
  agent
- |
  ageratum
- |
  Aggeus
- |
  aggie
- |
  agglomerate
- |
  agglutinate
- |
  agglutinated
- |
  aggrandize
- |
  aggrandizer
- |
  aggravate
- |
  aggravated
- |
  aggravating
- |
  aggravation
- |
  aggravator
- |
  aggregate
- |
  aggregation
- |
  aggregative
- |
  aggression
- |
  aggressive
- |
  aggressively
- |
  aggressor
- |
  aggrieve
- |
  aggrieved
- |
  aggrievedly
- |
  aggrievement
- |
  aghast
- |
  agile
- |
  agilely
- |
  agileness
- |
  agility
- |
  Agincourt
- |
  aging
- |
  agism
- |
  agist
- |
  agita
- |
  agitate
- |
  agitated
- |
  agitatedly
- |
  agitation
- |
  agitator
- |
  agitprop
- |
  agleam
- |
  aglitter
- |
  aglow
- |
  agnate
- |
  agnatic
- |
  agnation
- |
  Agnes
- |
  Agnew
- |
  agnostic
- |
  agnosticism
- |
  agonising
- |
  agonist
- |
  agonize
- |
  agonizing
- |
  agonizingly
- |
  agony
- |
  agora
- |
  agorae
- |
  agoraphobe
- |
  agoraphobia
- |
  agoraphobic
- |
  agrarian
- |
  agrarianism
- |
  agree
- |
  agreeable
- |
  agreeably
- |
  agreed
- |
  agreement
- |
  agribusiness
- |
  Agricola
- |
  agricultural
- |
  agriculture
- |
  Agrippa
- |
  Agrippina
- |
  agronomic
- |
  agronomical
- |
  agronomist
- |
  agronomy
- |
  aground
- |
  Aguinaldo
- |
  aguish
- |
  Agulhas
- |
  Ahaggar
- |
  ahead
- |
  ahimsa
- |
  Ahmadabad
- |
  Ahmedabad
- |
  aider
- |
  aigret
- |
  aigrette
- |
  Aiken
- |
  aikido
- |
  ailanthus
- |
  Aileen
- |
  aileron
- |
  ailing
- |
  ailment
- |
  aimless
- |
  aimlessly
- |
  aimlessness
- |
  aioli
- |
  airbag
- |
  airbase
- |
  airboat
- |
  airborne
- |
  airbrush
- |
  airbus
- |
  aircraft
- |
  airdrome
- |
  airdrop
- |
  Airedale
- |
  airfare
- |
  airfield
- |
  airflow
- |
  airfoil
- |
  airframe
- |
  airfreight
- |
  airhead
- |
  airily
- |
  airiness
- |
  airing
- |
  airless
- |
  airlessness
- |
  airlift
- |
  airline
- |
  airliner
- |
  airlock
- |
  airmail
- |
  airman
- |
  airmobile
- |
  airplane
- |
  airplay
- |
  airport
- |
  airpower
- |
  airship
- |
  airsick
- |
  airsickness
- |
  airspace
- |
  airstrike
- |
  airstrip
- |
  airtight
- |
  airtime
- |
  airwave
- |
  airwaves
- |
  airway
- |
  airwoman
- |
  airworthy
- |
  aisle
- |
  Aisne
- |
  aitch
- |
  Ajaccio
- |
  Akbar
- |
  Akhenaton
- |
  Akhmatova
- |
  Akhnaton
- |
  Akihito
- |
  akimbo
- |
  Akkad
- |
  Akkadian
- |
  Akron
- |
  akvavit
- |
  Alabama
- |
  Alabaman
- |
  Alabamian
- |
  alabaster
- |
  alacritous
- |
  alacrity
- |
  Aladdin
- |
  alameda
- |
  Alamo
- |
  Alamogordo
- |
  Alaric
- |
  alarm
- |
  alarmed
- |
  alarming
- |
  alarmingly
- |
  alarmism
- |
  alarmist
- |
  alarum
- |
  Alaska
- |
  Alaskan
- |
  albacore
- |
  Alban
- |
  Albania
- |
  Albanian
- |
  Albany
- |
  albatross
- |
  albedo
- |
  Albee
- |
  albeit
- |
  Albemarle
- |
  Albert
- |
  Alberta
- |
  Albertan
- |
  albescent
- |
  albinism
- |
  albino
- |
  Albion
- |
  Albireo
- |
  Alborg
- |
  Albright
- |
  album
- |
  albumen
- |
  albumin
- |
  albuminous
- |
  Albuquerque
- |
  alcaic
- |
  alcaics
- |
  alcalde
- |
  Alcatraz
- |
  alcazar
- |
  alchemic
- |
  alchemical
- |
  alchemically
- |
  alchemist
- |
  alchemize
- |
  alchemy
- |
  Alcibiades
- |
  alcohol
- |
  alcoholic
- |
  alcoholism
- |
  Alcor
- |
  Alcott
- |
  alcove
- |
  Alcuin
- |
  Alcyone
- |
  Aldabra
- |
  Aldan
- |
  Aldebaran
- |
  aldehyde
- |
  Alden
- |
  alder
- |
  alderman
- |
  Alderney
- |
  alderwoman
- |
  aleatoric
- |
  aleatory
- |
  alehouse
- |
  Alembert
- |
  alembic
- |
  Aleppo
- |
  alert
- |
  alertly
- |
  alertness
- |
  Aleut
- |
  Aleutian
- |
  Aleutians
- |
  alewife
- |
  alewives
- |
  Alexander
- |
  Alexandra
- |
  Alexandria
- |
  Alexandrian
- |
  alexandrine
- |
  alexia
- |
  Alexis
- |
  alfalfa
- |
  Alfonso
- |
  Alfred
- |
  Alfreda
- |
  alfresco
- |
  algae
- |
  algal
- |
  algebra
- |
  algebraic
- |
  Algenib
- |
  Alger
- |
  Algeria
- |
  Algerian
- |
  Algerine
- |
  Algernon
- |
  Algiers
- |
  Algol
- |
  Algonkian
- |
  Algonkin
- |
  Algonquian
- |
  Algonquin
- |
  algorithm
- |
  algorithmic
- |
  alias
- |
  alibi
- |
  Alicante
- |
  Alice
- |
  Alicia
- |
  alien
- |
  alienability
- |
  alienable
- |
  alienate
- |
  alienated
- |
  alienation
- |
  alienator
- |
  alienist
- |
  alienness
- |
  Alighieri
- |
  alight
- |
  align
- |
  aligner
- |
  alignment
- |
  alike
- |
  alikeness
- |
  aliment
- |
  alimentary
- |
  alimony
- |
  aline
- |
  alinement
- |
  Alioth
- |
  aliphatic
- |
  aliquot
- |
  Alison
- |
  Alistair
- |
  alive
- |
  aliveness
- |
  aliya
- |
  aliyah
- |
  alizarin
- |
  Alkaid
- |
  alkali
- |
  alkaline
- |
  alkalinity
- |
  alkalinize
- |
  alkalization
- |
  alkalize
- |
  alkaloid
- |
  alkaloidal
- |
  alkalosis
- |
  alkane
- |
  alkyd
- |
  Allah
- |
  Allahabad
- |
  Allan
- |
  allay
- |
  allee
- |
  allegation
- |
  allege
- |
  allegeable
- |
  alleged
- |
  allegedly
- |
  alleger
- |
  Alleghenies
- |
  Allegheny
- |
  allegiance
- |
  allegoric
- |
  allegorical
- |
  allegorist
- |
  allegorize
- |
  allegory
- |
  allegretto
- |
  allegro
- |
  allele
- |
  allelic
- |
  allelomorph
- |
  allelopathic
- |
  allelopathy
- |
  alleluia
- |
  Allen
- |
  Allende
- |
  Allentown
- |
  allergen
- |
  allergenic
- |
  allergic
- |
  allergically
- |
  allergist
- |
  allergy
- |
  alleviate
- |
  alleviation
- |
  alleviator
- |
  alley
- |
  alleyway
- |
  Allhallows
- |
  alliance
- |
  allied
- |
  alligator
- |
  Allison
- |
  alliterate
- |
  alliteration
- |
  alliterative
- |
  allocable
- |
  allocate
- |
  allocation
- |
  allocator
- |
  allocution
- |
  allomorph
- |
  allomorphic
- |
  allomorphism
- |
  allopathic
- |
  allopathist
- |
  allopathy
- |
  allophone
- |
  allophonic
- |
  allot
- |
  allotment
- |
  allotrope
- |
  allotropic
- |
  allotropical
- |
  allotropy
- |
  allotter
- |
  allover
- |
  allow
- |
  allowable
- |
  allowably
- |
  allowance
- |
  allowedly
- |
  alloy
- |
  allspice
- |
  allude
- |
  allure
- |
  allurement
- |
  alluring
- |
  alluringly
- |
  allusion
- |
  allusive
- |
  allusively
- |
  allusiveness
- |
  alluvia
- |
  alluvial
- |
  alluvion
- |
  alluvium
- |
  Allyn
- |
  Almach
- |
  almanac
- |
  almandite
- |
  Almaty
- |
  almightily
- |
  almightiness
- |
  Almighty
- |
  almighty
- |
  almond
- |
  almoner
- |
  almost
- |
  almsgiver
- |
  almshouse
- |
  aloes
- |
  aloft
- |
  aloha
- |
  alone
- |
  aloneness
- |
  along
- |
  alongshore
- |
  alongside
- |
  aloof
- |
  aloofly
- |
  aloofness
- |
  alopecia
- |
  aloud
- |
  Aloysius
- |
  alpaca
- |
  alpenhorn
- |
  alpha
- |
  alphabet
- |
  alphabetic
- |
  alphabetical
- |
  alphabetize
- |
  alphabetizer
- |
  alphameric
- |
  alphanumeric
- |
  Alphard
- |
  Alphecca
- |
  Alpheratz
- |
  Alphonso
- |
  Alpine
- |
  alpine
- |
  already
- |
  alright
- |
  Alsace
- |
  Alsatian
- |
  Altai
- |
  Altaic
- |
  Altair
- |
  altar
- |
  altarpiece
- |
  alter
- |
  alterable
- |
  alteration
- |
  altercate
- |
  altercation
- |
  alternate
- |
  alternately
- |
  alternation
- |
  alternative
- |
  alternator
- |
  Althea
- |
  altho
- |
  although
- |
  altimeter
- |
  altimetry
- |
  altiplano
- |
  altitude
- |
  altitudinal
- |
  altogether
- |
  Alton
- |
  Altoona
- |
  altruism
- |
  altruist
- |
  altruistic
- |
  alumina
- |
  aluminium
- |
  aluminize
- |
  aluminous
- |
  aluminum
- |
  alumna
- |
  alumnae
- |
  alumni
- |
  alumnus
- |
  Alvah
- |
  Alvarez
- |
  alveoli
- |
  alveolus
- |
  Alvin
- |
  always
- |
  Alyce
- |
  alyssum
- |
  Amagasaki
- |
  amain
- |
  amalgam
- |
  amalgamate
- |
  amalgamated
- |
  amalgamation
- |
  Amanda
- |
  amandine
- |
  amanuenses
- |
  amanuensis
- |
  amaranth
- |
  amaranthine
- |
  amaretto
- |
  Amarillo
- |
  amaryllis
- |
  amass
- |
  amasser
- |
  amassment
- |
  amateur
- |
  amateurish
- |
  amateurishly
- |
  amateurism
- |
  Amati
- |
  amative
- |
  amatively
- |
  amativeness
- |
  amatory
- |
  amaze
- |
  amazed
- |
  amazedly
- |
  amazement
- |
  amazing
- |
  amazingly
- |
  Amazon
- |
  amazon
- |
  Amazonia
- |
  Amazonian
- |
  amazonian
- |
  ambassador
- |
  ambassadress
- |
  Amber
- |
  amber
- |
  ambergris
- |
  ambiance
- |
  ambidextrous
- |
  ambience
- |
  ambient
- |
  ambiguity
- |
  ambiguous
- |
  ambiguously
- |
  ambit
- |
  ambition
- |
  ambitious
- |
  ambitiously
- |
  ambivalence
- |
  ambivalent
- |
  ambivalently
- |
  amble
- |
  ambler
- |
  Ambrose
- |
  ambrosia
- |
  ambrosial
- |
  ambulance
- |
  ambulant
- |
  ambulate
- |
  ambulation
- |
  ambulator
- |
  ambulatory
- |
  ambuscade
- |
  ambuscaded
- |
  ambuscader
- |
  ambush
- |
  ambusher
- |
  ameba
- |
  amebae
- |
  amebic
- |
  ameboid
- |
  Amelia
- |
  ameliorate
- |
  amelioration
- |
  ameliorative
- |
  ameliorator
- |
  amenability
- |
  amenable
- |
  amenableness
- |
  amenably
- |
  amend
- |
  amendable
- |
  amender
- |
  amendment
- |
  amends
- |
  Amenhotep
- |
  amenities
- |
  amenity
- |
  amenorrhea
- |
  amenorrheic
- |
  amenorrhoea
- |
  ament
- |
  Amerasian
- |
  amerce
- |
  amercement
- |
  America
- |
  American
- |
  Americana
- |
  Americanism
- |
  Americanize
- |
  Americanness
- |
  Americas
- |
  americium
- |
  Amerind
- |
  Amerindian
- |
  amethyst
- |
  amethystine
- |
  Amharic
- |
  Amherst
- |
  amiability
- |
  amiable
- |
  amiableness
- |
  amiably
- |
  amicability
- |
  amicable
- |
  amicably
- |
  amide
- |
  amidship
- |
  amidships
- |
  amidst
- |
  Amiens
- |
  amigo
- |
  amine
- |
  Amish
- |
  amiss
- |
  amity
- |
  Amman
- |
  ammeter
- |
  ammonia
- |
  ammonite
- |
  ammonium
- |
  ammunition
- |
  amnesia
- |
  amnesiac
- |
  amnesic
- |
  amnestic
- |
  amnesty
- |
  amnia
- |
  amnio
- |
  amnion
- |
  amnionic
- |
  amniotic
- |
  amoeba
- |
  amoebae
- |
  amoebic
- |
  amoeboid
- |
  among
- |
  amongst
- |
  amontillado
- |
  amoral
- |
  amoralism
- |
  amoralist
- |
  amorality
- |
  amorally
- |
  amorist
- |
  amorous
- |
  amorously
- |
  amorousness
- |
  amorphous
- |
  amorphously
- |
  amortizable
- |
  amortization
- |
  amortize
- |
  amount
- |
  amour
- |
  amoxicillin
- |
  amperage
- |
  Ampere
- |
  ampere
- |
  ampersand
- |
  amphetamine
- |
  amphibian
- |
  amphibious
- |
  amphibiously
- |
  amphibole
- |
  amphibolic
- |
  amphitheater
- |
  amphitheatre
- |
  amphora
- |
  amphorae
- |
  ampicillin
- |
  ample
- |
  ampleness
- |
  amplified
- |
  amplifier
- |
  amplify
- |
  amplitude
- |
  amply
- |
  ampoul
- |
  ampoule
- |
  ampul
- |
  ampule
- |
  ampulla
- |
  ampullae
- |
  amputate
- |
  amputation
- |
  amputator
- |
  amputee
- |
  Amritsar
- |
  Amsterdam
- |
  Amtrak
- |
  amuck
- |
  amulet
- |
  Amundsen
- |
  amusable
- |
  amuse
- |
  amused
- |
  amusedly
- |
  amusement
- |
  amusing
- |
  amusingly
- |
  amylase
- |
  Anabaptism
- |
  Anabaptist
- |
  anabolic
- |
  anabolism
- |
  anachronism
- |
  anachronous
- |
  anacolutha
- |
  anacoluthic
- |
  anacoluthon
- |
  anaconda
- |
  Anacreon
- |
  anaemia
- |
  anaemic
- |
  anaerobe
- |
  anaerobic
- |
  anaesthesia
- |
  anaesthetic
- |
  anaesthetist
- |
  anaesthetize
- |
  anagram
- |
  anagrammatic
- |
  Anaheim
- |
  analecta
- |
  analects
- |
  analgesia
- |
  analgesic
- |
  anally
- |
  analog
- |
  analogical
- |
  analogically
- |
  analogize
- |
  analogous
- |
  analogously
- |
  analogue
- |
  analogy
- |
  analysand
- |
  analyse
- |
  analyses
- |
  analysis
- |
  analyst
- |
  analytic
- |
  analytical
- |
  analytically
- |
  analyzable
- |
  analyze
- |
  analyzer
- |
  Ananias
- |
  anapaest
- |
  anapest
- |
  anapestic
- |
  anaphora
- |
  anaphoric
- |
  anarchic
- |
  anarchical
- |
  anarchically
- |
  anarchism
- |
  anarchist
- |
  anarchistic
- |
  anarchy
- |
  Anasazi
- |
  Anastasia
- |
  anastomoses
- |
  anastomosis
- |
  anathema
- |
  anathematize
- |
  Anatolia
- |
  Anatolian
- |
  anatomic
- |
  anatomical
- |
  anatomically
- |
  anatomist
- |
  anatomize
- |
  anatomy
- |
  Anaxagoras
- |
  ancestor
- |
  ancestral
- |
  ancestrally
- |
  ancestress
- |
  ancestry
- |
  anchor
- |
  Anchorage
- |
  anchorage
- |
  anchorite
- |
  anchoritic
- |
  anchorman
- |
  anchorperson
- |
  anchorwoman
- |
  anchovy
- |
  ancient
- |
  anciently
- |
  ancientness
- |
  ancients
- |
  ancillary
- |
  Andalusia
- |
  Andalusian
- |
  Andaman
- |
  Andamanese
- |
  andante
- |
  andantino
- |
  Andean
- |
  Andersen
- |
  Anderson
- |
  Andes
- |
  Andine
- |
  andiron
- |
  Andorra
- |
  Andorran
- |
  Andre
- |
  Andrea
- |
  Andrew
- |
  androgen
- |
  androgenic
- |
  androgyne
- |
  androgynous
- |
  androgyny
- |
  android
- |
  Andromeda
- |
  Andropov
- |
  Andros
- |
  anecdotal
- |
  anecdotalist
- |
  anecdotally
- |
  anecdote
- |
  anecdotist
- |
  anechoic
- |
  anemia
- |
  anemic
- |
  anemically
- |
  anemometer
- |
  anemone
- |
  anent
- |
  anerobic
- |
  aneroid
- |
  anesthesia
- |
  anesthetic
- |
  anesthetist
- |
  anesthetize
- |
  aneurism
- |
  aneurysm
- |
  aneurysmal
- |
  angel
- |
  Angela
- |
  Angeleno
- |
  angelfish
- |
  angelic
- |
  Angelica
- |
  angelica
- |
  angelical
- |
  angelically
- |
  Angelico
- |
  Angelina
- |
  Angeline
- |
  Angelo
- |
  Angelou
- |
  anger
- |
  Angers
- |
  angina
- |
  anginal
- |
  angiogenesis
- |
  angiogenic
- |
  angiogram
- |
  angiography
- |
  angioplasty
- |
  angiosperm
- |
  Angkor
- |
  Angle
- |
  angle
- |
  angled
- |
  angler
- |
  Angles
- |
  Anglesey
- |
  angleworm
- |
  Anglican
- |
  Anglicanism
- |
  Anglicism
- |
  Anglicize
- |
  anglicize
- |
  anglicized
- |
  angling
- |
  Anglo
- |
  Anglocentric
- |
  Anglophil
- |
  Anglophile
- |
  Anglophilia
- |
  Anglophobe
- |
  Anglophobia
- |
  Anglophobic
- |
  Anglophone
- |
  anglophone
- |
  Angola
- |
  Angolan
- |
  Angora
- |
  angora
- |
  angrily
- |
  angriness
- |
  angry
- |
  angst
- |
  angstrom
- |
  Anguilla
- |
  anguine
- |
  anguish
- |
  anguished
- |
  angular
- |
  angularity
- |
  angularly
- |
  Angus
- |
  anhydride
- |
  anhydrous
- |
  anilin
- |
  aniline
- |
  animadvert
- |
  animal
- |
  animalcule
- |
  animalism
- |
  animate
- |
  animated
- |
  animatedly
- |
  animation
- |
  animato
- |
  animator
- |
  anime
- |
  animism
- |
  animist
- |
  animistic
- |
  animosity
- |
  animus
- |
  anion
- |
  anionic
- |
  anionically
- |
  anise
- |
  aniseed
- |
  anisette
- |
  Anita
- |
  Anjou
- |
  Ankara
- |
  ankle
- |
  anklebone
- |
  anklet
- |
  ankylosis
- |
  ankylotic
- |
  Annabel
- |
  Annabelle
- |
  annalist
- |
  annalistic
- |
  annals
- |
  Annam
- |
  Annamese
- |
  Annapolis
- |
  Annapurna
- |
  anneal
- |
  annealer
- |
  annelid
- |
  Annenberg
- |
  Annetta
- |
  Annette
- |
  annex
- |
  annexation
- |
  annexe
- |
  annexed
- |
  Annie
- |
  annihilate
- |
  annihilation
- |
  annihilator
- |
  anniversary
- |
  annotate
- |
  annotation
- |
  annotative
- |
  annotator
- |
  announce
- |
  announcement
- |
  announcer
- |
  annoy
- |
  annoyance
- |
  annoyed
- |
  annoying
- |
  annoyingly
- |
  annual
- |
  annually
- |
  annuitant
- |
  annuity
- |
  annul
- |
  annular
- |
  annularity
- |
  annularly
- |
  annuli
- |
  annulment
- |
  annulus
- |
  annunciate
- |
  Annunciation
- |
  annunciation
- |
  annunciator
- |
  anodal
- |
  anode
- |
  anodic
- |
  anodize
- |
  anodyne
- |
  anoint
- |
  anointed
- |
  anointer
- |
  anointment
- |
  anole
- |
  anomalistic
- |
  anomalous
- |
  anomalously
- |
  anomaly
- |
  anomie
- |
  anomy
- |
  anonymity
- |
  anonymous
- |
  anonymously
- |
  anopheles
- |
  anorak
- |
  anorectic
- |
  anorexia
- |
  anorexic
- |
  another
- |
  Anouilh
- |
  Anselm
- |
  Anshan
- |
  answer
- |
  answerable
- |
  answerably
- |
  answerer
- |
  antacid
- |
  antagonise
- |
  antagonism
- |
  antagonist
- |
  antagonistic
- |
  antagonize
- |
  Antalya
- |
  Antananarivo
- |
  Antarctic
- |
  antarctic
- |
  Antarctica
- |
  Antares
- |
  anteater
- |
  antebellum
- |
  antecede
- |
  antecedence
- |
  antecedent
- |
  antecedents
- |
  antechamber
- |
  antedate
- |
  antediluvian
- |
  antelope
- |
  antenna
- |
  antennae
- |
  antepenult
- |
  anterior
- |
  anteriority
- |
  anteriorly
- |
  anteroom
- |
  anthem
- |
  anther
- |
  anthill
- |
  anthologist
- |
  anthologize
- |
  anthology
- |
  Anthony
- |
  anthracite
- |
  anthracitic
- |
  anthrax
- |
  anthropoid
- |
  anthropology
- |
  antiabortion
- |
  antiaging
- |
  antiaircraft
- |
  antialcohol
- |
  antiallergic
- |
  antianxiety
- |
  antibiotic
- |
  antibody
- |
  antic
- |
  anticancer
- |
  Antichrist
- |
  antichrist
- |
  anticipate
- |
  anticipation
- |
  anticipator
- |
  anticipatory
- |
  anticlerical
- |
  anticlimax
- |
  anticline
- |
  anticolonial
- |
  anticrime
- |
  antics
- |
  anticyclone
- |
  anticyclonic
- |
  antidotal
- |
  antidote
- |
  antidrug
- |
  Antietam
- |
  antifascism
- |
  antifascist
- |
  antifeminism
- |
  antifeminist
- |
  antifreeze
- |
  antifungal
- |
  antigen
- |
  antigenic
- |
  antigenicity
- |
  Antigone
- |
  antigravity
- |
  Antigua
- |
  Antiguan
- |
  antihero
- |
  antiheroic
- |
  antiheroine
- |
  antihumanism
- |
  antiknock
- |
  antilabor
- |
  antiliberal
- |
  Antillean
- |
  Antilles
- |
  antilock
- |
  antilog
- |
  antimacassar
- |
  antimalarial
- |
  antimatter
- |
  antimissile
- |
  antimitotic
- |
  antimonial
- |
  antimonic
- |
  antimonous
- |
  antimony
- |
  antinarcotic
- |
  antinausea
- |
  antineutron
- |
  antinoise
- |
  antinomian
- |
  antinomy
- |
  antinovel
- |
  antinuclear
- |
  Antioch
- |
  antioxidant
- |
  antipacifist
- |
  antiparticle
- |
  antipasti
- |
  antipasto
- |
  antipathetic
- |
  antipathy
- |
  antiphon
- |
  antiphonal
- |
  antiphonally
- |
  antiphony
- |
  antipodal
- |
  antipode
- |
  antipodean
- |
  Antipodes
- |
  antipodes
- |
  antipole
- |
  antipope
- |
  antipoverty
- |
  antiproton
- |
  antipyresis
- |
  antipyretic
- |
  antiquarian
- |
  antiquary
- |
  antiquate
- |
  antiquated
- |
  antiquation
- |
  antique
- |
  antiquely
- |
  antiqueness
- |
  antiquer
- |
  antiquities
- |
  antiquity
- |
  antiradical
- |
  antirational
- |
  antis
- |
  antisemite
- |
  antisemitic
- |
  antisemitism
- |
  antisepsis
- |
  antiseptic
- |
  antisera
- |
  antiserum
- |
  antislavery
- |
  antismoking
- |
  antisocial
- |
  antisocially
- |
  antistatic
- |
  antistrophe
- |
  antitakeover
- |
  antitank
- |
  antitheft
- |
  antitheses
- |
  antithesis
- |
  antithetic
- |
  antithetical
- |
  antitoxic
- |
  antitoxin
- |
  antitrust
- |
  antitumor
- |
  antitussive
- |
  antiunion
- |
  antivenin
- |
  antiviral
- |
  antivirus
- |
  antiwar
- |
  antler
- |
  antlered
- |
  Antlia
- |
  Antoinette
- |
  Anton
- |
  Antonia
- |
  Antonio
- |
  Antonius
- |
  Antony
- |
  antonym
- |
  antonymic
- |
  antonymous
- |
  antonymy
- |
  Antrim
- |
  antsy
- |
  Antwerp
- |
  Anubis
- |
  anvil
- |
  anxiety
- |
  anxious
- |
  anxiously
- |
  anxiousness
- |
  anybody
- |
  anyhow
- |
  anymore
- |
  anyone
- |
  anyplace
- |
  anything
- |
  anytime
- |
  anyway
- |
  anywhere
- |
  anywise
- |
  Aorangi
- |
  aorist
- |
  aoristic
- |
  aorta
- |
  aortae
- |
  aortal
- |
  aortic
- |
  aoudad
- |
  apace
- |
  Apache
- |
  Apachean
- |
  apanage
- |
  apart
- |
  apartheid
- |
  apartment
- |
  apartness
- |
  apathetic
- |
  apathy
- |
  apatite
- |
  apatosaur
- |
  apatosaurus
- |
  apelike
- |
  Apennine
- |
  Apennines
- |
  apercu
- |
  aperitif
- |
  apertural
- |
  aperture
- |
  aphasia
- |
  aphasiac
- |
  aphasic
- |
  aphelia
- |
  aphelian
- |
  aphelion
- |
  apheresis
- |
  aphid
- |
  aphides
- |
  aphis
- |
  aphorism
- |
  aphorist
- |
  aphoristic
- |
  aphorize
- |
  aphrodisiac
- |
  Aphrodite
- |
  apiarian
- |
  apiarist
- |
  apiary
- |
  apical
- |
  apically
- |
  apices
- |
  apicultural
- |
  apiculture
- |
  apiculturist
- |
  apiece
- |
  aplenty
- |
  aplomb
- |
  apnea
- |
  Apocalypse
- |
  apocalypse
- |
  apocalyptic
- |
  Apocrypha
- |
  apocrypha
- |
  Apocryphal
- |
  apocryphal
- |
  apocryphally
- |
  apodeictic
- |
  apodictic
- |
  apogee
- |
  apolitical
- |
  apolitically
- |
  Apollo
- |
  apollo
- |
  Apollonian
- |
  Apollonius
- |
  apologetic
- |
  apologetical
- |
  apologetics
- |
  apologia
- |
  apologise
- |
  apologist
- |
  apologize
- |
  apologue
- |
  apology
- |
  apophthegm
- |
  apoplectic
- |
  apoplexy
- |
  aporia
- |
  aport
- |
  apostasy
- |
  apostate
- |
  apostatical
- |
  apostatize
- |
  Apostle
- |
  apostle
- |
  apostleship
- |
  apostolic
- |
  apostrophe
- |
  apostrophic
- |
  apostrophize
- |
  apothecary
- |
  apothegm
- |
  apothegmatic
- |
  apothem
- |
  apotheoses
- |
  apotheosis
- |
  apotheosize
- |
  appal
- |
  Appalachia
- |
  Appalachian
- |
  Appalachians
- |
  appall
- |
  appalled
- |
  appalling
- |
  appallingly
- |
  Appaloosa
- |
  appaloosa
- |
  appanage
- |
  apparatchik
- |
  apparatchiki
- |
  apparatus
- |
  apparel
- |
  apparent
- |
  apparently
- |
  apparition
- |
  apparitional
- |
  appeal
- |
  appealable
- |
  appealer
- |
  appealing
- |
  appealingly
- |
  appear
- |
  appearance
- |
  appeasable
- |
  appease
- |
  appeasement
- |
  appeaser
- |
  appellant
- |
  appellate
- |
  appellation
- |
  appellee
- |
  append
- |
  appendage
- |
  appendectomy
- |
  appendices
- |
  appendicitis
- |
  appendix
- |
  appertain
- |
  appetency
- |
  appetite
- |
  appetitive
- |
  appetizer
- |
  appetizing
- |
  appetizingly
- |
  applaud
- |
  applaudable
- |
  applauder
- |
  applause
- |
  apple
- |
  applejack
- |
  applesauce
- |
  applet
- |
  Appleton
- |
  appliance
- |
  applicable
- |
  applicably
- |
  applicant
- |
  application
- |
  applications
- |
  applicator
- |
  applied
- |
  applier
- |
  applique
- |
  appliqued
- |
  apply
- |
  appoint
- |
  appointed
- |
  appointee
- |
  appointive
- |
  appointment
- |
  appointments
- |
  Appomattox
- |
  apportion
- |
  appose
- |
  apposite
- |
  appositely
- |
  appositeness
- |
  apposition
- |
  appositional
- |
  appositive
- |
  appraisable
- |
  appraisal
- |
  appraise
- |
  appraisement
- |
  appraiser
- |
  appraisingly
- |
  appreciable
- |
  appreciably
- |
  appreciate
- |
  appreciation
- |
  appreciative
- |
  appreciator
- |
  appreciatory
- |
  apprehend
- |
  apprehension
- |
  apprehensive
- |
  apprentice
- |
  apprise
- |
  apprize
- |
  approach
- |
  approachable
- |
  approbation
- |
  approbative
- |
  approbatory
- |
  appropriate
- |
  appropriator
- |
  approval
- |
  approve
- |
  approvingly
- |
  approximate
- |
  appurtenance
- |
  appurtenant
- |
  apricot
- |
  April
- |
  apriorism
- |
  apron
- |
  aproned
- |
  apropos
- |
  apsidal
- |
  apsides
- |
  apsis
- |
  aptitude
- |
  aptly
- |
  aptness
- |
  Apuleius
- |
  Aqaba
- |
  aquaculture
- |
  aquae
- |
  aquamarine
- |
  aquanaut
- |
  aquaplane
- |
  aquaplaning
- |
  aquaria
- |
  Aquarian
- |
  aquarium
- |
  Aquarius
- |
  aquatic
- |
  aquatically
- |
  aquatics
- |
  aquatint
- |
  aquavit
- |
  aqueduct
- |
  aqueous
- |
  aquiculture
- |
  aquifer
- |
  Aquila
- |
  aquiline
- |
  Aquinas
- |
  Aquino
- |
  Aquitaine
- |
  Arabella
- |
  arabesque
- |
  Arabia
- |
  Arabian
- |
  Arabic
- |
  arability
- |
  arable
- |
  arachnid
- |
  arachnidan
- |
  Arafat
- |
  Arafura
- |
  Aragon
- |
  Aragonese
- |
  Araguaia
- |
  Araguaya
- |
  Aramaic
- |
  aramid
- |
  Arapaho
- |
  Arapahoe
- |
  Ararat
- |
  Arawak
- |
  Arawakan
- |
  Arbela
- |
  Arbil
- |
  arbiter
- |
  arbitrage
- |
  arbitrager
- |
  arbitrageur
- |
  arbitrament
- |
  arbitrarily
- |
  arbitrary
- |
  arbitrate
- |
  arbitration
- |
  arbitrator
- |
  arbor
- |
  arboreal
- |
  arboreta
- |
  arboretum
- |
  arborvitae
- |
  arbour
- |
  arbovirus
- |
  arbutus
- |
  arcade
- |
  arcaded
- |
  Arcadia
- |
  Arcadian
- |
  arcading
- |
  Arcady
- |
  arcana
- |
  arcane
- |
  arcanum
- |
  archaeologic
- |
  archaeology
- |
  archaic
- |
  archaically
- |
  archaism
- |
  archaist
- |
  archaistic
- |
  Archangel
- |
  archangel
- |
  archbishop
- |
  archdeacon
- |
  archdeaconry
- |
  archdiocesan
- |
  archdiocese
- |
  archduchess
- |
  archduchy
- |
  archduke
- |
  Archean
- |
  arched
- |
  archenemy
- |
  archeology
- |
  Archeozoic
- |
  archer
- |
  archerfish
- |
  archery
- |
  archetypal
- |
  archetype
- |
  archetypic
- |
  archetypical
- |
  Archfiend
- |
  archfiend
- |
  Archibald
- |
  Archie
- |
  Archimedean
- |
  Archimedes
- |
  archipelagic
- |
  archipelago
- |
  architect
- |
  architecture
- |
  architrave
- |
  archival
- |
  archive
- |
  archives
- |
  archivist
- |
  archly
- |
  archness
- |
  archon
- |
  archrival
- |
  archway
- |
  Arctic
- |
  arctic
- |
  Arcturus
- |
  arcuate
- |
  Ardabil
- |
  Ardebil
- |
  Ardell
- |
  Ardelle
- |
  Arden
- |
  ardency
- |
  Ardennes
- |
  ardent
- |
  ardently
- |
  ardor
- |
  ardour
- |
  arduous
- |
  arduously
- |
  arduousness
- |
  areal
- |
  areaway
- |
  arena
- |
  areola
- |
  areolae
- |
  areolar
- |
  areolate
- |
  Arequipa
- |
  arete
- |
  argent
- |
  Argentina
- |
  Argentine
- |
  Argentinean
- |
  Argentinian
- |
  argentite
- |
  Argolis
- |
  argon
- |
  Argonaut
- |
  argonaut
- |
  Argonne
- |
  Argos
- |
  argosy
- |
  argot
- |
  arguable
- |
  arguably
- |
  argue
- |
  arguer
- |
  argument
- |
  argumentive
- |
  Argus
- |
  argyle
- |
  argyll
- |
  Arhus
- |
  aridity
- |
  aridly
- |
  aridness
- |
  Aries
- |
  aright
- |
  Ariosto
- |
  arise
- |
  arisen
- |
  Aristides
- |
  aristocracy
- |
  aristocrat
- |
  aristocratic
- |
  Aristophanes
- |
  Aristotelian
- |
  Aristotle
- |
  arithmetic
- |
  arithmetical
- |
  Arius
- |
  Arizona
- |
  Arizonan
- |
  Arizonian
- |
  Arkansan
- |
  Arkansas
- |
  Arkhangelsk
- |
  Arkwright
- |
  Arleen
- |
  Arlen
- |
  Arlene
- |
  Arlin
- |
  Arline
- |
  Arlington
- |
  armada
- |
  armadillo
- |
  Armageddon
- |
  Armagh
- |
  armament
- |
  armaments
- |
  Armand
- |
  armature
- |
  armband
- |
  armchair
- |
  armed
- |
  Armenia
- |
  Armenian
- |
  armful
- |
  armhole
- |
  armistice
- |
  armless
- |
  armlet
- |
  armoire
- |
  armor
- |
  armored
- |
  armorer
- |
  armorial
- |
  armory
- |
  armour
- |
  armoured
- |
  armoury
- |
  armpit
- |
  armrest
- |
  armsful
- |
  Armstrong
- |
  armyworm
- |
  Arnhem
- |
  arnica
- |
  Arnold
- |
  aroma
- |
  aromatherapy
- |
  aromatic
- |
  aromatically
- |
  aromaticity
- |
  aromatics
- |
  arose
- |
  around
- |
  arousal
- |
  arouse
- |
  aroused
- |
  arousing
- |
  Arpanet
- |
  arpeggiate
- |
  arpeggiation
- |
  arpeggio
- |
  arraign
- |
  arraignment
- |
  arrange
- |
  arrangement
- |
  arranger
- |
  arrant
- |
  arras
- |
  array
- |
  arrear
- |
  arrearage
- |
  arrears
- |
  arrest
- |
  arrester
- |
  arresting
- |
  arrestor
- |
  arrhythmia
- |
  arrhythmic
- |
  arrhythmical
- |
  arrival
- |
  arrive
- |
  arrivederci
- |
  arriviste
- |
  arrogance
- |
  arrogant
- |
  arrogantly
- |
  arrogate
- |
  arrogation
- |
  arrogative
- |
  arrow
- |
  arrowhead
- |
  arrowroot
- |
  arroyo
- |
  arsenal
- |
  arsenic
- |
  arsenical
- |
  arson
- |
  arsonist
- |
  Artaxerxes
- |
  artefact
- |
  Artemis
- |
  arterial
- |
  arteriolar
- |
  arteriole
- |
  artery
- |
  artesian
- |
  artful
- |
  artfully
- |
  artfulness
- |
  arthritic
- |
  arthritides
- |
  arthritis
- |
  arthropod
- |
  arthroscope
- |
  arthroscopic
- |
  arthroscopy
- |
  Arthur
- |
  Arthurian
- |
  artichoke
- |
  article
- |
  articulable
- |
  articulacy
- |
  articular
- |
  articulate
- |
  articulately
- |
  articulation
- |
  articulator
- |
  artifact
- |
  artifactual
- |
  artifice
- |
  artificer
- |
  artificial
- |
  artificially
- |
  artillerist
- |
  artillery
- |
  artilleryman
- |
  artily
- |
  artiness
- |
  artisan
- |
  artisanal
- |
  artisanship
- |
  artist
- |
  artiste
- |
  artistic
- |
  artistically
- |
  artistry
- |
  artless
- |
  artlessly
- |
  artlessness
- |
  artsy
- |
  artwork
- |
  Aruba
- |
  arugula
- |
  Aryan
- |
  asafetida
- |
  asafoetida
- |
  Asama
- |
  asbestos
- |
  asbestosis
- |
  ascend
- |
  ascendancy
- |
  ascendant
- |
  ascendency
- |
  ascendent
- |
  Ascension
- |
  ascension
- |
  ascent
- |
  ascertain
- |
  ascesis
- |
  ascetic
- |
  ascetically
- |
  asceticism
- |
  ASCII
- |
  Asclepius
- |
  ascot
- |
  ascribable
- |
  ascribe
- |
  ascription
- |
  asepsis
- |
  aseptic
- |
  asexual
- |
  asexuality
- |
  asexually
- |
  ashamed
- |
  ashamedly
- |
  Ashanti
- |
  ashcan
- |
  ashen
- |
  ashes
- |
  Ashgabat
- |
  Ashkenazi
- |
  Ashkenazic
- |
  Ashkenazim
- |
  Ashkhabad
- |
  ashlar
- |
  Ashley
- |
  ashore
- |
  ashram
- |
  ashtray
- |
  Asian
- |
  Asiatic
- |
  aside
- |
  Asimov
- |
  asinine
- |
  asininely
- |
  asininity
- |
  askance
- |
  asker
- |
  askew
- |
  aslant
- |
  asleep
- |
  Asmara
- |
  Asmera
- |
  asocial
- |
  asparagus
- |
  aspartame
- |
  aspect
- |
  aspen
- |
  asperities
- |
  asperity
- |
  asperse
- |
  aspersion
- |
  aspersions
- |
  asphalt
- |
  asphaltic
- |
  asphaltum
- |
  asphodel
- |
  asphyxia
- |
  asphyxiate
- |
  asphyxiation
- |
  asphyxiator
- |
  aspic
- |
  aspidistra
- |
  aspirant
- |
  aspirate
- |
  aspiration
- |
  aspirational
- |
  aspirations
- |
  aspirator
- |
  aspire
- |
  aspirer
- |
  aspirin
- |
  aspiring
- |
  aspiringly
- |
  asquint
- |
  Asquith
- |
  Assad
- |
  assail
- |
  assailable
- |
  assailant
- |
  assailer
- |
  assassin
- |
  assassinate
- |
  assault
- |
  assaulter
- |
  assaultive
- |
  assay
- |
  assayable
- |
  assayer
- |
  assemblage
- |
  assemble
- |
  assembler
- |
  Assembly
- |
  assembly
- |
  assemblyman
- |
  assent
- |
  assenter
- |
  assentor
- |
  assert
- |
  asserter
- |
  assertion
- |
  assertive
- |
  assertively
- |
  assertor
- |
  assess
- |
  assessable
- |
  assessment
- |
  assessor
- |
  asset
- |
  assets
- |
  asseverate
- |
  asseveration
- |
  asshole
- |
  assiduities
- |
  assiduity
- |
  assiduous
- |
  assiduously
- |
  assign
- |
  assignable
- |
  assignation
- |
  assignee
- |
  assigner
- |
  assignment
- |
  assignor
- |
  assimilable
- |
  assimilate
- |
  assimilation
- |
  assimilative
- |
  assimilator
- |
  assimilatory
- |
  Assiniboin
- |
  assist
- |
  assistance
- |
  assistant
- |
  assize
- |
  assizes
- |
  associate
- |
  associated
- |
  association
- |
  associative
- |
  assonance
- |
  assonant
- |
  assonantal
- |
  assonate
- |
  assort
- |
  assortative
- |
  assorted
- |
  assorter
- |
  assortment
- |
  assuage
- |
  assuagement
- |
  assumable
- |
  assumably
- |
  assume
- |
  assumed
- |
  assumedly
- |
  assuming
- |
  Assumption
- |
  assumption
- |
  assumptive
- |
  assurance
- |
  assure
- |
  assured
- |
  assuredly
- |
  assuredness
- |
  assurer
- |
  assuror
- |
  Assyria
- |
  Assyrian
- |
  Astaire
- |
  astatine
- |
  aster
- |
  asterisk
- |
  astern
- |
  asteroid
- |
  asthma
- |
  asthmatic
- |
  astigmatic
- |
  astigmatism
- |
  astir
- |
  astonish
- |
  astonished
- |
  astonishing
- |
  astonishment
- |
  Astor
- |
  astound
- |
  astounded
- |
  astounding
- |
  astoundingly
- |
  astraddle
- |
  Astrakhan
- |
  astrakhan
- |
  astral
- |
  astray
- |
  Astrid
- |
  astride
- |
  astringency
- |
  astringent
- |
  astringently
- |
  astrobiology
- |
  astrolabe
- |
  astrologer
- |
  astrologic
- |
  astrological
- |
  astrologist
- |
  astrology
- |
  astronaut
- |
  astronautic
- |
  astronautics
- |
  astronomer
- |
  astronomic
- |
  astronomical
- |
  astronomy
- |
  astrophysics
- |
  AstroTurf
- |
  Asturias
- |
  astute
- |
  astutely
- |
  astuteness
- |
  Asuncion
- |
  asunder
- |
  Aswan
- |
  asylum
- |
  asymmetric
- |
  asymmetrical
- |
  asymmetry
- |
  asymptomatic
- |
  asymptote
- |
  asymptotic
- |
  asymptotical
- |
  Asyut
- |
  Atacama
- |
  ataractic
- |
  ataraxia
- |
  ataraxic
- |
  ataraxy
- |
  Ataturk
- |
  atavism
- |
  atavist
- |
  atavistic
- |
  ataxia
- |
  ataxic
- |
  Atchafalaya
- |
  atelier
- |
  Athabasca
- |
  Athabascan
- |
  Athabaska
- |
  Athabaskan
- |
  Athapaskan
- |
  atheism
- |
  atheist
- |
  atheistic
- |
  atheistical
- |
  Athena
- |
  athenaeum
- |
  Athene
- |
  atheneum
- |
  Athenian
- |
  Athens
- |
  athirst
- |
  athlete
- |
  athletic
- |
  athletically
- |
  athleticism
- |
  athletics
- |
  athwart
- |
  atilt
- |
  Atlanta
- |
  Atlantan
- |
  Atlantic
- |
  Atlantis
- |
  Atlas
- |
  atlas
- |
  atlatl
- |
  Atman
- |
  atman
- |
  atmosphere
- |
  atmospheric
- |
  atmospherics
- |
  atoll
- |
  atomic
- |
  atomically
- |
  atomism
- |
  atomist
- |
  atomistic
- |
  atomization
- |
  atomize
- |
  atomizer
- |
  atonal
- |
  atonalism
- |
  atonalist
- |
  atonality
- |
  atonally
- |
  atone
- |
  atonement
- |
  atoner
- |
  atria
- |
  atrial
- |
  atrium
- |
  atrocious
- |
  atrociously
- |
  atrocity
- |
  atrophic
- |
  atrophied
- |
  atrophy
- |
  atropin
- |
  atropine
- |
  Atropos
- |
  attach
- |
  attachable
- |
  attache
- |
  attached
- |
  attachment
- |
  attack
- |
  attacker
- |
  attacking
- |
  attain
- |
  attainable
- |
  attainder
- |
  attainment
- |
  attaint
- |
  attar
- |
  attempt
- |
  attemptable
- |
  attempted
- |
  Attenborough
- |
  attend
- |
  attendance
- |
  attendant
- |
  attendee
- |
  attention
- |
  attentions
- |
  attentive
- |
  attentively
- |
  attenuate
- |
  attenuated
- |
  attenuation
- |
  attest
- |
  attestation
- |
  attester
- |
  attestor
- |
  Attic
- |
  attic
- |
  Attica
- |
  Atticism
- |
  atticism
- |
  Attila
- |
  attire
- |
  attitude
- |
  attitudinal
- |
  attitudinize
- |
  Attlee
- |
  attorney
- |
  attorneyship
- |
  attract
- |
  attractable
- |
  attractant
- |
  attracted
- |
  attraction
- |
  attractive
- |
  attractively
- |
  attributable
- |
  attribute
- |
  attributer
- |
  attribution
- |
  attributive
- |
  attributor
- |
  attrit
- |
  attrition
- |
  attritional
- |
  Attucks
- |
  attune
- |
  attuned
- |
  attunement
- |
  atwitter
- |
  Atwood
- |
  atypical
- |
  atypically
- |
  aubergine
- |
  Aubrey
- |
  auburn
- |
  Auckland
- |
  auction
- |
  auctioneer
- |
  auctorial
- |
  audacious
- |
  audaciously
- |
  audacity
- |
  Auden
- |
  audial
- |
  audibility
- |
  audible
- |
  audibly
- |
  audience
- |
  audio
- |
  audiobook
- |
  audiological
- |
  audiologist
- |
  audiology
- |
  audiometer
- |
  audiometric
- |
  audiophile
- |
  audiotape
- |
  audiovisual
- |
  audiovisuals
- |
  audit
- |
  audition
- |
  auditor
- |
  auditoria
- |
  auditorium
- |
  auditory
- |
  Audra
- |
  Audrey
- |
  Audubon
- |
  auger
- |
  aught
- |
  augment
- |
  augmentation
- |
  augmentative
- |
  augmenter
- |
  Augsburg
- |
  augur
- |
  augural
- |
  augury
- |
  August
- |
  august
- |
  Augusta
- |
  Augustan
- |
  Augustine
- |
  Augustinian
- |
  augustly
- |
  augustness
- |
  Augustus
- |
  aurae
- |
  aural
- |
  aurally
- |
  Aurangabad
- |
  aurar
- |
  aureate
- |
  Aurelia
- |
  Aurelian
- |
  Aurelius
- |
  aureola
- |
  aureole
- |
  auricle
- |
  auricled
- |
  auricular
- |
  Aurora
- |
  aurora
- |
  aurorae
- |
  auroral
- |
  Aurungabad
- |
  Auschwitz
- |
  auscultate
- |
  auscultation
- |
  auspice
- |
  auspices
- |
  auspicious
- |
  auspiciously
- |
  Aussie
- |
  Austen
- |
  austere
- |
  austerely
- |
  austerity
- |
  Austerlitz
- |
  Austin
- |
  Austral
- |
  austral
- |
  Australasia
- |
  Australasian
- |
  Australia
- |
  Australian
- |
  Australoid
- |
  Austria
- |
  Austrian
- |
  Austronesia
- |
  Austronesian
- |
  autarch
- |
  autarchic
- |
  autarchy
- |
  autarkic
- |
  autarky
- |
  auteur
- |
  auteurism
- |
  auteurist
- |
  authentic
- |
  authenticate
- |
  authenticity
- |
  author
- |
  authoress
- |
  authorial
- |
  authorise
- |
  authorities
- |
  authority
- |
  authorize
- |
  authorship
- |
  autism
- |
  autistic
- |
  autobahn
- |
  autochthon
- |
  autochthones
- |
  autoclave
- |
  autocracy
- |
  autocrat
- |
  autocratic
- |
  autocratical
- |
  autodidact
- |
  autodidactic
- |
  autograph
- |
  autographic
- |
  autoimmune
- |
  autoimmunity
- |
  automata
- |
  automate
- |
  automated
- |
  automatic
- |
  automation
- |
  automatism
- |
  automatize
- |
  automaton
- |
  automobile
- |
  automotive
- |
  autonomic
- |
  autonomist
- |
  autonomous
- |
  autonomously
- |
  autonomy
- |
  autopilot
- |
  autopsied
- |
  autopsist
- |
  autopsy
- |
  autosome
- |
  autotroph
- |
  autotrophic
- |
  autoworker
- |
  autumn
- |
  autumnal
- |
  Auvergne
- |
  auxiliaries
- |
  auxiliary
- |
  auxin
- |
  avail
- |
  availability
- |
  available
- |
  avalanche
- |
  avarice
- |
  avaricious
- |
  avariciously
- |
  avast
- |
  avatar
- |
  avaunt
- |
  avenge
- |
  avenger
- |
  avenue
- |
  average
- |
  averagely
- |
  averment
- |
  averral
- |
  Averroes
- |
  averse
- |
  aversely
- |
  aversion
- |
  aversive
- |
  avert
- |
  avertable
- |
  avertible
- |
  avian
- |
  aviarist
- |
  aviary
- |
  aviation
- |
  aviator
- |
  aviatrices
- |
  aviatrix
- |
  Avicenna
- |
  avidity
- |
  avidly
- |
  avidness
- |
  Avignon
- |
  avionic
- |
  avionics
- |
  avitaminosis
- |
  avocado
- |
  avocation
- |
  avocational
- |
  avocet
- |
  avoid
- |
  avoidable
- |
  avoidably
- |
  avoidance
- |
  avoider
- |
  avoirdupois
- |
  avouch
- |
  avowal
- |
  avowed
- |
  avowedly
- |
  avuncular
- |
  AWACS
- |
  await
- |
  awake
- |
  awaken
- |
  awakening
- |
  award
- |
  aware
- |
  awareness
- |
  awash
- |
  aweigh
- |
  awesome
- |
  awesomely
- |
  awesomeness
- |
  awestricken
- |
  awestruck
- |
  awful
- |
  awfully
- |
  awfulness
- |
  awhile
- |
  awhirl
- |
  awkward
- |
  awkwardly
- |
  awkwardness
- |
  awned
- |
  awning
- |
  awoke
- |
  awoken
- |
  axial
- |
  axially
- |
  axilla
- |
  axillae
- |
  axiom
- |
  axiomatic
- |
  axletree
- |
  Axminster
- |
  axolotl
- |
  ayatollah
- |
  Aylesbury
- |
  Aymara
- |
  Aymaran
- |
  Ayrshire
- |
  azalea
- |
  Azcapotzalco
- |
  Azerbaijan
- |
  Azerbaijani
- |
  azimuth
- |
  azimuthal
- |
  Azorean
- |
  Azores
- |
  Azorian
- |
  Aztec
- |
  Aztecan
- |
  azure
- |
  Baalim
- |
  Babar
- |
  Babbitt
- |
  babbitt
- |
  Babbittry
- |
  babble
- |
  babbler
- |
  Babel
- |
  babel
- |
  Baber
- |
  Babette
- |
  Babism
- |
  baboon
- |
  Babur
- |
  babushka
- |
  babyhood
- |
  babyish
- |
  Babylon
- |
  Babylonia
- |
  Babylonian
- |
  babysat
- |
  babysit
- |
  babysitter
- |
  babysitting
- |
  babytalk
- |
  Bacall
- |
  baccarat
- |
  bacchanal
- |
  Bacchanalia
- |
  bacchanalia
- |
  Bacchanalian
- |
  bacchanalian
- |
  Bacchic
- |
  Bacchus
- |
  bachelor
- |
  bachelordom
- |
  bachelorette
- |
  bachelorhood
- |
  bacillar
- |
  bacillary
- |
  bacilli
- |
  bacillus
- |
  bacitracin
- |
  backache
- |
  backbeat
- |
  backbench
- |
  backbencher
- |
  backbit
- |
  backbite
- |
  backbiter
- |
  backbiting
- |
  backbitten
- |
  backboard
- |
  backbone
- |
  backbreaking
- |
  backcourt
- |
  backdate
- |
  backdoor
- |
  backdrop
- |
  backer
- |
  backfield
- |
  backfire
- |
  backgammon
- |
  background
- |
  backgrounder
- |
  backhand
- |
  backhanded
- |
  backhandedly
- |
  backhoe
- |
  backing
- |
  backlash
- |
  backless
- |
  backlight
- |
  backlog
- |
  backpack
- |
  backpacker
- |
  backpacking
- |
  backpedal
- |
  backrest
- |
  backroom
- |
  backseat
- |
  backsheesh
- |
  backside
- |
  backslap
- |
  backslapper
- |
  backslapping
- |
  backslash
- |
  backslid
- |
  backslidden
- |
  backslide
- |
  backslider
- |
  backspace
- |
  backspin
- |
  backstage
- |
  backstair
- |
  backstairs
- |
  backstop
- |
  backstretch
- |
  backstroke
- |
  backswept
- |
  backswing
- |
  backtalk
- |
  backtrack
- |
  backup
- |
  backward
- |
  backwardly
- |
  backwardness
- |
  backwards
- |
  backwash
- |
  backwater
- |
  backwoods
- |
  backwoodsman
- |
  backyard
- |
  Bacon
- |
  bacon
- |
  bacteria
- |
  bacterial
- |
  bacterially
- |
  bactericidal
- |
  bactericide
- |
  bacteriology
- |
  bacterium
- |
  Bactria
- |
  Bactrian
- |
  Baden
- |
  badge
- |
  badger
- |
  badinage
- |
  badland
- |
  Badlands
- |
  badlands
- |
  badly
- |
  badman
- |
  badminton
- |
  badmouth
- |
  badness
- |
  Baedeker
- |
  Baffin
- |
  baffle
- |
  baffled
- |
  bafflement
- |
  baffler
- |
  baffling
- |
  bagasse
- |
  bagatelle
- |
  Bagdad
- |
  bagel
- |
  bagful
- |
  baggage
- |
  bagger
- |
  Baggie
- |
  baggie
- |
  Baggies
- |
  baggily
- |
  bagginess
- |
  baggy
- |
  Baghdad
- |
  bagman
- |
  bagnio
- |
  bagpipe
- |
  bagpiper
- |
  bagpipes
- |
  baguette
- |
  Baguio
- |
  Bahai
- |
  Bahaman
- |
  Bahamanian
- |
  Bahamas
- |
  Bahamian
- |
  Bahia
- |
  Bahrain
- |
  Bahraini
- |
  Bahrein
- |
  Baikal
- |
  bailable
- |
  bailee
- |
  bailer
- |
  Bailey
- |
  bailiff
- |
  bailiwick
- |
  bailor
- |
  bailout
- |
  bailsman
- |
  Bairiki
- |
  bairn
- |
  baiter
- |
  baiza
- |
  baize
- |
  Bakelite
- |
  Baker
- |
  baker
- |
  Bakersfield
- |
  bakery
- |
  bakeshop
- |
  Bakhtaran
- |
  baking
- |
  baklava
- |
  baksheesh
- |
  Bakunin
- |
  balaclava
- |
  balalaika
- |
  balance
- |
  balanced
- |
  Balanchine
- |
  Balaton
- |
  Balboa
- |
  balboa
- |
  balbriggan
- |
  balcony
- |
  baldachin
- |
  baldachino
- |
  balderdash
- |
  baldfaced
- |
  balding
- |
  baldly
- |
  baldness
- |
  baldric
- |
  Baldwin
- |
  baleen
- |
  baleful
- |
  balefully
- |
  balefulness
- |
  baler
- |
  Balfour
- |
  Balikpapan
- |
  Balinese
- |
  Balkan
- |
  Balkans
- |
  balker
- |
  Balkhash
- |
  balky
- |
  ballad
- |
  ballade
- |
  balladeer
- |
  balladry
- |
  ballast
- |
  ballboy
- |
  ballcarrier
- |
  ballcock
- |
  ballerina
- |
  ballet
- |
  balletic
- |
  balletomane
- |
  ballgame
- |
  ballgirl
- |
  ballistic
- |
  ballistics
- |
  balloon
- |
  balloonist
- |
  ballot
- |
  balloter
- |
  balloting
- |
  ballpark
- |
  ballplayer
- |
  ballpoint
- |
  ballroom
- |
  balls
- |
  ballute
- |
  Ballycastle
- |
  ballyhoo
- |
  Ballymena
- |
  Ballymoney
- |
  ballyrag
- |
  balmily
- |
  balminess
- |
  balmy
- |
  baloney
- |
  balsa
- |
  balsam
- |
  balsamic
- |
  Baltic
- |
  Baltimore
- |
  baluster
- |
  balustrade
- |
  balustraded
- |
  Balzac
- |
  Bamako
- |
  bamboo
- |
  bamboozle
- |
  banal
- |
  banality
- |
  banally
- |
  banana
- |
  Banaras
- |
  Banares
- |
  Banbridge
- |
  bandage
- |
  bandaid
- |
  bandana
- |
  bandanna
- |
  bandbox
- |
  bandeau
- |
  bandeaux
- |
  banded
- |
  bander
- |
  banderol
- |
  banderole
- |
  bandicoot
- |
  bandit
- |
  banditry
- |
  bandmaster
- |
  bandoleer
- |
  bandolier
- |
  bandsaw
- |
  bandsman
- |
  bandstand
- |
  Bandung
- |
  bandwagon
- |
  bandwidth
- |
  bandy
- |
  bandylegged
- |
  baneful
- |
  Bangalore
- |
  Bangkok
- |
  Bangladesh
- |
  Bangladeshi
- |
  bangle
- |
  Bangor
- |
  bangs
- |
  Bangui
- |
  banian
- |
  banish
- |
  banishment
- |
  banister
- |
  Banjermasin
- |
  banjo
- |
  banjoist
- |
  Banjul
- |
  bankable
- |
  bankbook
- |
  bankcard
- |
  banker
- |
  banking
- |
  banknote
- |
  bankroll
- |
  bankrupt
- |
  bankruptcy
- |
  banks
- |
  Banneker
- |
  banner
- |
  banning
- |
  Bannister
- |
  bannister
- |
  bannock
- |
  banns
- |
  banquet
- |
  banqueter
- |
  banquette
- |
  banshee
- |
  banshie
- |
  bantam
- |
  bantamweight
- |
  banter
- |
  bantering
- |
  banteringly
- |
  Bantu
- |
  Bantustan
- |
  banyan
- |
  banzai
- |
  baobab
- |
  Baotou
- |
  baptism
- |
  baptismal
- |
  Baptist
- |
  baptist
- |
  baptistery
- |
  baptistry
- |
  baptize
- |
  baptizer
- |
  Barabbas
- |
  Barbadian
- |
  Barbados
- |
  Barbara
- |
  barbarian
- |
  barbarianism
- |
  barbaric
- |
  barbarism
- |
  barbarity
- |
  barbarize
- |
  Barbarossa
- |
  barbarous
- |
  barbarously
- |
  Barbary
- |
  barbecue
- |
  barbed
- |
  barbel
- |
  barbell
- |
  barbeque
- |
  barber
- |
  barberry
- |
  barbershop
- |
  barbital
- |
  barbiturate
- |
  Barbuda
- |
  Barbudan
- |
  barbwire
- |
  barcarole
- |
  barcarolle
- |
  Barcelona
- |
  Barclay
- |
  bardic
- |
  bareback
- |
  barebacked
- |
  barefaced
- |
  barefacedly
- |
  barefoot
- |
  barefooted
- |
  barehanded
- |
  bareheaded
- |
  Bareilly
- |
  barelegged
- |
  barely
- |
  bareness
- |
  barfly
- |
  bargain
- |
  bargainer
- |
  bargaining
- |
  barge
- |
  bargeman
- |
  barite
- |
  baritone
- |
  barium
- |
  barkeep
- |
  barkeeper
- |
  barker
- |
  Barking
- |
  barley
- |
  barmaid
- |
  barman
- |
  Barnabas
- |
  Barnaby
- |
  barnacle
- |
  barnacled
- |
  Barnard
- |
  Barnaul
- |
  Barnet
- |
  Barnett
- |
  Barney
- |
  barnstorm
- |
  barnstormer
- |
  Barnum
- |
  barnyard
- |
  Baroda
- |
  barograph
- |
  barographic
- |
  barometer
- |
  barometric
- |
  barometrical
- |
  barometry
- |
  baron
- |
  baronage
- |
  baroness
- |
  baronet
- |
  baronetcy
- |
  baronetess
- |
  baronial
- |
  barony
- |
  Baroque
- |
  baroque
- |
  baroquely
- |
  barouche
- |
  barque
- |
  Barquisimeto
- |
  barrack
- |
  barracking
- |
  barracks
- |
  barracuda
- |
  barrage
- |
  Barranquilla
- |
  barratry
- |
  barre
- |
  barred
- |
  barrel
- |
  barreled
- |
  barrelhead
- |
  barren
- |
  barrenness
- |
  barrens
- |
  Barrett
- |
  barrette
- |
  barricade
- |
  Barrie
- |
  barrier
- |
  barring
- |
  barrio
- |
  barrister
- |
  barroom
- |
  barrow
- |
  Barry
- |
  Barrymore
- |
  bartender
- |
  barter
- |
  barterer
- |
  Barth
- |
  Barthes
- |
  Bartholdi
- |
  Bartholomew
- |
  Bartlett
- |
  Bartok
- |
  Barton
- |
  Baruch
- |
  baryon
- |
  Baryshnikov
- |
  basal
- |
  basally
- |
  basalt
- |
  basaltic
- |
  baseball
- |
  baseboard
- |
  baseborn
- |
  based
- |
  Basel
- |
  baseless
- |
  baselessness
- |
  baseline
- |
  basely
- |
  baseman
- |
  basement
- |
  baseness
- |
  basenji
- |
  bases
- |
  basher
- |
  bashful
- |
  bashfully
- |
  bashfulness
- |
  bashing
- |
  BASIC
- |
  Basic
- |
  basic
- |
  basically
- |
  basicity
- |
  basics
- |
  Basie
- |
  Basil
- |
  basil
- |
  Basilan
- |
  Basildon
- |
  basilica
- |
  basilican
- |
  basilisk
- |
  basin
- |
  basinal
- |
  basinful
- |
  basis
- |
  basket
- |
  basketball
- |
  basketful
- |
  basketry
- |
  basketwork
- |
  Basle
- |
  Basque
- |
  Basra
- |
  basset
- |
  Basseterre
- |
  bassi
- |
  bassinet
- |
  bassist
- |
  basso
- |
  bassoon
- |
  bassoonist
- |
  basswood
- |
  bastard
- |
  bastardize
- |
  bastardly
- |
  bastardy
- |
  baste
- |
  baster
- |
  bastile
- |
  Bastille
- |
  bastille
- |
  bastinade
- |
  bastinado
- |
  bastion
- |
  bastioned
- |
  Basutoland
- |
  Bataan
- |
  Batavia
- |
  batch
- |
  bateau
- |
  bateaux
- |
  bated
- |
  bathe
- |
  bather
- |
  bathetic
- |
  bathhouse
- |
  bathing
- |
  bathmat
- |
  bathos
- |
  bathrobe
- |
  bathroom
- |
  baths
- |
  Bathsheba
- |
  bathtub
- |
  Bathurst
- |
  bathyscaph
- |
  bathyscaphe
- |
  bathysphere
- |
  batik
- |
  Batista
- |
  batiste
- |
  Batman
- |
  batman
- |
  baton
- |
  batsman
- |
  battalion
- |
  batten
- |
  batter
- |
  battered
- |
  batterer
- |
  battering
- |
  battery
- |
  batting
- |
  battle
- |
  battleax
- |
  battleaxe
- |
  battledore
- |
  battlefield
- |
  battlefront
- |
  battleground
- |
  battlement
- |
  battlemented
- |
  battlements
- |
  battler
- |
  battleship
- |
  battlewagon
- |
  batty
- |
  bauble
- |
  Baudelaire
- |
  Baudouin
- |
  Bauhaus
- |
  baulk
- |
  bauxite
- |
  Bavaria
- |
  Bavarian
- |
  bawdily
- |
  bawdiness
- |
  bawdy
- |
  bawdyhouse
- |
  bawler
- |
  Bayamon
- |
  bayberry
- |
  Baykal
- |
  bayonet
- |
  bayou
- |
  Bayreuth
- |
  bazaar
- |
  bazar
- |
  bazooka
- |
  beach
- |
  beachcomber
- |
  beachcombing
- |
  beachhead
- |
  beacon
- |
  beading
- |
  beadle
- |
  beads
- |
  beady
- |
  beagle
- |
  beaked
- |
  beaker
- |
  beanbag
- |
  beanball
- |
  beanie
- |
  beano
- |
  beanpole
- |
  bearable
- |
  bearably
- |
  beard
- |
  bearded
- |
  beardless
- |
  Beardsley
- |
  bearer
- |
  bearing
- |
  bearings
- |
  bearish
- |
  bearishly
- |
  bearishness
- |
  bearlike
- |
  bearskin
- |
  beast
- |
  beastliness
- |
  beastly
- |
  beatable
- |
  beaten
- |
  beater
- |
  beatific
- |
  beatifically
- |
  beatify
- |
  beating
- |
  beatitude
- |
  Beatitudes
- |
  Beatles
- |
  beatnik
- |
  Beatrice
- |
  Beatrix
- |
  Beaufort
- |
  Beauharnais
- |
  Beaujolais
- |
  Beaumarchais
- |
  Beaumont
- |
  Beauregard
- |
  beaut
- |
  beauteous
- |
  beauteously
- |
  beautician
- |
  beautifier
- |
  beautiful
- |
  beautifully
- |
  beautify
- |
  beauty
- |
  Beauvoir
- |
  beaux
- |
  beaver
- |
  beaverboard
- |
  Beaverton
- |
  bebop
- |
  becalm
- |
  became
- |
  because
- |
  bechamel
- |
  Bechuana
- |
  Bechuanaland
- |
  Becket
- |
  Beckett
- |
  beckon
- |
  Becky
- |
  becloud
- |
  become
- |
  becoming
- |
  becomingly
- |
  bedaub
- |
  bedazzle
- |
  bedazzlement
- |
  bedbug
- |
  bedclothes
- |
  bedcover
- |
  bedding
- |
  bedeck
- |
  bedevil
- |
  bedevilment
- |
  bedew
- |
  bedfast
- |
  bedfellow
- |
  Bedford
- |
  Bedfordshire
- |
  bedim
- |
  bedizen
- |
  bedlam
- |
  bedlinen
- |
  Bedloe
- |
  Bedouin
- |
  bedouin
- |
  bedpan
- |
  bedpost
- |
  bedraggle
- |
  bedraggled
- |
  bedridden
- |
  bedrock
- |
  bedroll
- |
  bedroom
- |
  bedside
- |
  bedsore
- |
  bedspread
- |
  bedstead
- |
  bedtime
- |
  Beduin
- |
  beduin
- |
  bedwetting
- |
  beech
- |
  beechen
- |
  Beecher
- |
  beechnut
- |
  beefalo
- |
  beefburger
- |
  beefcake
- |
  beefeater
- |
  beefiness
- |
  beefsteak
- |
  beefy
- |
  beehive
- |
  beekeeper
- |
  beekeeping
- |
  beeline
- |
  Beelzebub
- |
  beeper
- |
  Beerbohm
- |
  Beersheba
- |
  beery
- |
  beeswax
- |
  Beethoven
- |
  beetle
- |
  Beeton
- |
  beetroot
- |
  beeves
- |
  befall
- |
  befallen
- |
  befell
- |
  befit
- |
  befitting
- |
  befog
- |
  before
- |
  beforehand
- |
  befoul
- |
  befriend
- |
  befuddle
- |
  befuddled
- |
  befuddlement
- |
  began
- |
  begat
- |
  beget
- |
  begetter
- |
  beggar
- |
  beggarliness
- |
  beggarly
- |
  beggary
- |
  Begin
- |
  begin
- |
  beginner
- |
  beginning
- |
  beginnings
- |
  begone
- |
  begonia
- |
  begot
- |
  begotten
- |
  begrime
- |
  begrudge
- |
  begrudgingly
- |
  beguile
- |
  beguilement
- |
  beguiler
- |
  beguiling
- |
  beguilingly
- |
  beguine
- |
  begum
- |
  begun
- |
  behalf
- |
  Behan
- |
  behave
- |
  behavior
- |
  behavioral
- |
  behaviorism
- |
  behaviorist
- |
  behaviour
- |
  behavioural
- |
  behead
- |
  beheld
- |
  behemoth
- |
  behest
- |
  behind
- |
  behindhand
- |
  behold
- |
  beholden
- |
  beholder
- |
  behoof
- |
  behoove
- |
  beige
- |
  Beijing
- |
  being
- |
  Beira
- |
  Beirut
- |
  bejewel
- |
  bejeweled
- |
  bejewelled
- |
  belabor
- |
  belabour
- |
  Belarus
- |
  belated
- |
  belatedly
- |
  belatedness
- |
  Belau
- |
  belay
- |
  belch
- |
  beldam
- |
  beldame
- |
  beleaguer
- |
  beleaguered
- |
  Belem
- |
  Belfast
- |
  belfry
- |
  Belgian
- |
  Belgium
- |
  Belgorod
- |
  Belgrade
- |
  belie
- |
  belief
- |
  believable
- |
  believably
- |
  believe
- |
  believer
- |
  belike
- |
  Belinda
- |
  belittle
- |
  belittlement
- |
  belittler
- |
  Belize
- |
  Belizean
- |
  Bella
- |
  belladonna
- |
  Bellatrix
- |
  bellbottom
- |
  bellbottomed
- |
  bellboy
- |
  Belle
- |
  belle
- |
  belletrism
- |
  belletrist
- |
  belletristic
- |
  Bellevue
- |
  bellflower
- |
  bellhop
- |
  bellicose
- |
  bellicosity
- |
  belligerence
- |
  belligerency
- |
  belligerent
- |
  Bellini
- |
  bellman
- |
  Bellow
- |
  bellow
- |
  bellows
- |
  bellwether
- |
  belly
- |
  bellyache
- |
  bellybutton
- |
  bellyful
- |
  Belmopan
- |
  belong
- |
  belonging
- |
  belongings
- |
  Belorussia
- |
  Belorussian
- |
  beloved
- |
  below
- |
  belowdecks
- |
  Belshazzar
- |
  Beltway
- |
  beltway
- |
  beluga
- |
  belvedere
- |
  bemire
- |
  bemoan
- |
  bemuse
- |
  bemused
- |
  bemusedly
- |
  bemusement
- |
  Benares
- |
  Bench
- |
  bench
- |
  benchmark
- |
  benchwarmer
- |
  bendable
- |
  bender
- |
  bends
- |
  beneath
- |
  Benedict
- |
  Benedictine
- |
  Benediction
- |
  benediction
- |
  benedictory
- |
  benefaction
- |
  benefactor
- |
  benefactress
- |
  benefice
- |
  beneficed
- |
  beneficence
- |
  beneficent
- |
  beneficently
- |
  beneficial
- |
  beneficially
- |
  beneficiary
- |
  benefit
- |
  Benelux
- |
  Benet
- |
  benevolence
- |
  benevolent
- |
  benevolently
- |
  Bengal
- |
  Bengalese
- |
  Bengali
- |
  Benghazi
- |
  benighted
- |
  benightedly
- |
  benign
- |
  benignancy
- |
  benignant
- |
  benignantly
- |
  benignity
- |
  benignly
- |
  Benin
- |
  Beninese
- |
  benison
- |
  Benjamin
- |
  Bennett
- |
  Bennie
- |
  Benny
- |
  Bentham
- |
  benthic
- |
  Benton
- |
  bentonite
- |
  bentwood
- |
  benumb
- |
  Benxi
- |
  Benzedrine
- |
  benzene
- |
  benzine
- |
  benzoate
- |
  benzocaine
- |
  benzoin
- |
  benzol
- |
  Beograd
- |
  Beowulf
- |
  bequeath
- |
  bequeathal
- |
  bequeather
- |
  bequeathment
- |
  bequest
- |
  berate
- |
  Berber
- |
  berceuse
- |
  bereave
- |
  bereaved
- |
  bereavement
- |
  bereft
- |
  Berenice
- |
  beret
- |
  Bergen
- |
  Bergman
- |
  Bergson
- |
  beriberi
- |
  Bering
- |
  Berkeley
- |
  Berkeleyite
- |
  berkelium
- |
  Berkshire
- |
  Berkshires
- |
  Berlin
- |
  Berliner
- |
  Berlioz
- |
  Bermuda
- |
  Bermudan
- |
  Bermudas
- |
  bermudas
- |
  Bermudian
- |
  Bernadette
- |
  Bernadine
- |
  Bernard
- |
  Berne
- |
  Bernese
- |
  Bernhard
- |
  Bernhardt
- |
  Bernice
- |
  Bernie
- |
  Bernini
- |
  Bernstein
- |
  Berra
- |
  Berry
- |
  berry
- |
  berrylike
- |
  berserk
- |
  berth
- |
  Bertha
- |
  berthed
- |
  Bertram
- |
  Bertrand
- |
  Beryl
- |
  beryl
- |
  berylline
- |
  beryllium
- |
  beseech
- |
  beseecher
- |
  beseeching
- |
  beseechingly
- |
  beseem
- |
  beset
- |
  besetting
- |
  beside
- |
  besides
- |
  besiege
- |
  besieger
- |
  Beskids
- |
  besmear
- |
  besmirch
- |
  besmircher
- |
  besom
- |
  besot
- |
  besotted
- |
  besought
- |
  bespangle
- |
  bespatter
- |
  bespeak
- |
  bespoke
- |
  bespoken
- |
  besprinkle
- |
  Bessarabia
- |
  Bessarabian
- |
  Bessemer
- |
  Bessie
- |
  bestial
- |
  bestiality
- |
  bestialize
- |
  bestially
- |
  bestiary
- |
  bestir
- |
  bestow
- |
  bestowal
- |
  bestrew
- |
  bestrewn
- |
  bestrid
- |
  bestridden
- |
  bestride
- |
  bestrode
- |
  bestseller
- |
  bestselling
- |
  betake
- |
  betaken
- |
  betatron
- |
  betcha
- |
  betel
- |
  Betelgeuse
- |
  bethel
- |
  Bethesda
- |
  bethink
- |
  Bethlehem
- |
  bethought
- |
  Bethune
- |
  betide
- |
  betimes
- |
  Betjeman
- |
  betoken
- |
  betook
- |
  betray
- |
  betrayal
- |
  betrayer
- |
  betroth
- |
  betrothal
- |
  betrothed
- |
  Betsey
- |
  Betsy
- |
  betta
- |
  Bette
- |
  better
- |
  betterment
- |
  betters
- |
  Bettie
- |
  betting
- |
  bettor
- |
  Betty
- |
  Bettye
- |
  between
- |
  betwixt
- |
  Beulah
- |
  bevel
- |
  beveled
- |
  beverage
- |
  Beverley
- |
  Beverly
- |
  bewail
- |
  beware
- |
  bewigged
- |
  bewilder
- |
  bewildered
- |
  bewildering
- |
  bewilderment
- |
  bewitch
- |
  bewitched
- |
  bewitching
- |
  bewitchingly
- |
  bewitchment
- |
  Bexley
- |
  beyond
- |
  bezel
- |
  bhang
- |
  Bharat
- |
  Bhopal
- |
  Bhutan
- |
  Bhutanese
- |
  Bhutto
- |
  Biafra
- |
  Biafran
- |
  Bialystok
- |
  biannual
- |
  biannually
- |
  Biarritz
- |
  biased
- |
  biathlon
- |
  bibelot
- |
  Bible
- |
  bible
- |
  Biblical
- |
  biblical
- |
  Biblically
- |
  bibliography
- |
  bibliophile
- |
  bibliophilic
- |
  bibliophily
- |
  bibulous
- |
  bibulously
- |
  bicameral
- |
  bicameralism
- |
  bicarb
- |
  bicarbonate
- |
  bicentenary
- |
  bicentennial
- |
  biceps
- |
  bicker
- |
  bickerer
- |
  bickering
- |
  biconcave
- |
  biconcavity
- |
  biconvex
- |
  biconvexity
- |
  bicuspid
- |
  bicycle
- |
  bicycler
- |
  bicyclist
- |
  biddable
- |
  bidden
- |
  bidder
- |
  bidding
- |
  biddy
- |
  bidet
- |
  Bielefeld
- |
  biennia
- |
  biennial
- |
  biennially
- |
  biennium
- |
  Bierce
- |
  bifocal
- |
  bifocals
- |
  bifurcate
- |
  bifurcation
- |
  bigamist
- |
  bigamous
- |
  bigamy
- |
  Bigfoot
- |
  bigfoot
- |
  biggie
- |
  biggish
- |
  bighearted
- |
  bighorn
- |
  bight
- |
  bigmouth
- |
  bigness
- |
  bigot
- |
  bigoted
- |
  bigotry
- |
  bigshot
- |
  bigwig
- |
  bijou
- |
  bijoux
- |
  biker
- |
  bikeway
- |
  Bikini
- |
  bikini
- |
  bilateral
- |
  bilaterality
- |
  bilaterally
- |
  Bilbao
- |
  bilge
- |
  biliary
- |
  bilingual
- |
  bilingualism
- |
  bilingually
- |
  bilious
- |
  biliously
- |
  biliousness
- |
  bilker
- |
  billable
- |
  billboard
- |
  billed
- |
  billet
- |
  billfold
- |
  billiard
- |
  billiards
- |
  Billie
- |
  billing
- |
  Billings
- |
  billingsgate
- |
  billion
- |
  billionaire
- |
  billionth
- |
  billow
- |
  billowy
- |
  Billy
- |
  billy
- |
  Biloxi
- |
  bimbo
- |
  bimetal
- |
  bimetallic
- |
  bimetallism
- |
  Biminis
- |
  bimodal
- |
  bimodality
- |
  bimonthly
- |
  binary
- |
  binational
- |
  binaural
- |
  binaurally
- |
  binder
- |
  bindery
- |
  binding
- |
  binge
- |
  binger
- |
  Bingham
- |
  bingo
- |
  binnacle
- |
  binocular
- |
  binocularly
- |
  binoculars
- |
  binomial
- |
  binomially
- |
  biochemical
- |
  biochemist
- |
  biochemistry
- |
  biodegrade
- |
  biodiversity
- |
  bioengineer
- |
  bioethical
- |
  bioethicist
- |
  bioethics
- |
  biofeedback
- |
  biogas
- |
  biogenesis
- |
  biogenetic
- |
  biogenic
- |
  biogeography
- |
  biographer
- |
  biographic
- |
  biographical
- |
  biography
- |
  Bioko
- |
  biologic
- |
  biological
- |
  biologically
- |
  biologist
- |
  biology
- |
  biomass
- |
  biome
- |
  biomechanics
- |
  biomedical
- |
  biomedicine
- |
  bionic
- |
  bionically
- |
  bionics
- |
  biophysical
- |
  biophysicist
- |
  biophysics
- |
  biopic
- |
  biopsy
- |
  bioreserve
- |
  biorhythm
- |
  biorhythmic
- |
  biosphere
- |
  biospheric
- |
  biosynthesis
- |
  biosynthetic
- |
  biota
- |
  biotech
- |
  biotic
- |
  biotin
- |
  biotite
- |
  bipartisan
- |
  bipartite
- |
  biped
- |
  bipedal
- |
  biplane
- |
  bipolar
- |
  bipolarity
- |
  biracial
- |
  biracialism
- |
  birch
- |
  birchen
- |
  birdbath
- |
  birdbrain
- |
  birdbrained
- |
  birder
- |
  birdhouse
- |
  birdie
- |
  birding
- |
  birdlime
- |
  birdseed
- |
  birdshot
- |
  birdwatcher
- |
  birdwatching
- |
  biretta
- |
  Birkenhead
- |
  Birmingham
- |
  birth
- |
  birthday
- |
  birthmark
- |
  birthplace
- |
  birthrate
- |
  birthright
- |
  birthstone
- |
  Bisayas
- |
  Biscay
- |
  biscuit
- |
  bisect
- |
  bisection
- |
  bisector
- |
  bisexual
- |
  bisexualism
- |
  bisexuality
- |
  bisexually
- |
  Bishkek
- |
  bishop
- |
  bishopric
- |
  Bismarck
- |
  Bismarckian
- |
  bismuth
- |
  bison
- |
  bisque
- |
  Bissau
- |
  bistro
- |
  bitch
- |
  bitchily
- |
  bitchiness
- |
  bitchy
- |
  biter
- |
  bitewing
- |
  Bithynia
- |
  Bithynian
- |
  biting
- |
  bitingly
- |
  bitten
- |
  bitter
- |
  bitterly
- |
  bittern
- |
  bitterness
- |
  bitters
- |
  bittersweet
- |
  bittiness
- |
  bitty
- |
  bitumen
- |
  bituminous
- |
  bivalent
- |
  bivalve
- |
  bivouac
- |
  biweekly
- |
  biyearly
- |
  bizarre
- |
  bizarrely
- |
  bizarreness
- |
  bizarrerie
- |
  Bizet
- |
  blabber
- |
  blabbermouth
- |
  Black
- |
  black
- |
  blackamoor
- |
  blackball
- |
  blackberry
- |
  blackbird
- |
  blackboard
- |
  blackbody
- |
  Blackburn
- |
  blackcurrant
- |
  blacken
- |
  blackened
- |
  blackener
- |
  blackface
- |
  Blackfeet
- |
  blackfish
- |
  Blackfoot
- |
  blackguard
- |
  blackguardly
- |
  blackhead
- |
  blacking
- |
  blackish
- |
  blackjack
- |
  blacklight
- |
  blacklist
- |
  blackly
- |
  blackmail
- |
  blackmailer
- |
  Blackmun
- |
  blackness
- |
  blackout
- |
  Blackpool
- |
  blacksmith
- |
  blacksnake
- |
  Blackstone
- |
  blackthorn
- |
  blacktop
- |
  Blackwell
- |
  bladder
- |
  blade
- |
  bladed
- |
  blading
- |
  blain
- |
  Blaine
- |
  Blair
- |
  Blake
- |
  blamable
- |
  blamably
- |
  blame
- |
  blameable
- |
  blameless
- |
  blamelessly
- |
  blameworthy
- |
  Blanc
- |
  Blanch
- |
  blanch
- |
  Blanche
- |
  blancmange
- |
  bland
- |
  blandish
- |
  blandisher
- |
  blandishment
- |
  blandly
- |
  blandness
- |
  blank
- |
  blanket
- |
  blankly
- |
  blankness
- |
  blanquette
- |
  Blantyre
- |
  blare
- |
  blarney
- |
  blase
- |
  blaspheme
- |
  blasphemer
- |
  blasphemous
- |
  blasphemy
- |
  blast
- |
  blasted
- |
  blaster
- |
  blasting
- |
  blastoff
- |
  blatancy
- |
  blatant
- |
  blatantly
- |
  blather
- |
  blatherer
- |
  blatherskite
- |
  blaze
- |
  blazer
- |
  blazes
- |
  blazing
- |
  blazon
- |
  blazonry
- |
  bleach
- |
  bleacher
- |
  bleachers
- |
  bleak
- |
  bleakish
- |
  bleakly
- |
  bleakness
- |
  blear
- |
  blearily
- |
  bleariness
- |
  bleary
- |
  bleat
- |
  bleed
- |
  bleeder
- |
  bleeding
- |
  bleep
- |
  blemish
- |
  blemished
- |
  blench
- |
  blend
- |
  blender
- |
  blent
- |
  bless
- |
  blessed
- |
  blessedly
- |
  blessedness
- |
  blessing
- |
  blest
- |
  blether
- |
  Bligh
- |
  blight
- |
  blighted
- |
  blimp
- |
  blind
- |
  blinder
- |
  blinders
- |
  blindfold
- |
  blindfolded
- |
  blinding
- |
  blindingly
- |
  blindly
- |
  blindness
- |
  blindside
- |
  blink
- |
  blinker
- |
  blinkers
- |
  blintz
- |
  blintze
- |
  bliss
- |
  blissful
- |
  blissfully
- |
  blissfulness
- |
  blister
- |
  blistered
- |
  blistering
- |
  blisteringly
- |
  blistery
- |
  blithe
- |
  blitheful
- |
  blithefully
- |
  blithely
- |
  blitheness
- |
  blither
- |
  blithesome
- |
  blithesomely
- |
  blitz
- |
  blitzkrieg
- |
  blizzard
- |
  bloat
- |
  bloated
- |
  block
- |
  blockade
- |
  blockader
- |
  blockage
- |
  blockbuster
- |
  blockbusting
- |
  blocker
- |
  blockhead
- |
  blockhouse
- |
  Bloemfontein
- |
  bloke
- |
  blond
- |
  blonde
- |
  blondish
- |
  blondness
- |
  blood
- |
  bloodbath
- |
  blooded
- |
  bloodhound
- |
  bloodily
- |
  bloodiness
- |
  bloodless
- |
  bloodlessly
- |
  bloodletting
- |
  bloodline
- |
  bloodmobile
- |
  bloodroot
- |
  bloodshed
- |
  bloodshot
- |
  bloodstain
- |
  bloodstained
- |
  bloodstock
- |
  bloodstream
- |
  bloodsucker
- |
  bloodsucking
- |
  bloodthirsty
- |
  bloody
- |
  bloom
- |
  Bloomer
- |
  bloomer
- |
  bloomers
- |
  Bloomfield
- |
  blooming
- |
  Bloomington
- |
  bloomy
- |
  blooper
- |
  blossom
- |
  blossoming
- |
  blossomy
- |
  blotch
- |
  blotched
- |
  blotchiness
- |
  blotchy
- |
  blotter
- |
  blouse
- |
  blower
- |
  blowfly
- |
  blowgun
- |
  blowhard
- |
  blowhole
- |
  blown
- |
  blowout
- |
  blowpipe
- |
  blowsy
- |
  blowtorch
- |
  blowup
- |
  blowy
- |
  blowzy
- |
  blubber
- |
  blubbery
- |
  bludgeon
- |
  Bluebeard
- |
  bluebell
- |
  blueberry
- |
  bluebird
- |
  blueblood
- |
  bluebonnet
- |
  bluebottle
- |
  bluefish
- |
  bluegill
- |
  bluegrass
- |
  blueing
- |
  blueish
- |
  bluejacket
- |
  bluejay
- |
  bluejeans
- |
  blueness
- |
  Bluenose
- |
  bluenose
- |
  bluenosed
- |
  bluepoint
- |
  blueprint
- |
  blues
- |
  bluesman
- |
  bluestocking
- |
  bluesy
- |
  bluet
- |
  bluets
- |
  bluff
- |
  bluffer
- |
  bluffly
- |
  bluffness
- |
  bluing
- |
  bluish
- |
  blunder
- |
  blunderbuss
- |
  blunderer
- |
  blunderingly
- |
  blunt
- |
  bluntly
- |
  bluntness
- |
  blurb
- |
  blurred
- |
  blurriness
- |
  blurry
- |
  blurt
- |
  blush
- |
  blusher
- |
  blushful
- |
  bluster
- |
  blusterer
- |
  blustery
- |
  Boadicea
- |
  board
- |
  boarder
- |
  boardroom
- |
  boards
- |
  boardwalk
- |
  boast
- |
  boaster
- |
  boastful
- |
  boastfully
- |
  boastfulness
- |
  boatel
- |
  boater
- |
  boathouse
- |
  boating
- |
  boatman
- |
  boatswain
- |
  Bobbie
- |
  bobbin
- |
  bobble
- |
  Bobby
- |
  bobby
- |
  bobbysocks
- |
  bobbysox
- |
  bobbysoxer
- |
  bobcat
- |
  bobolink
- |
  bobsled
- |
  bobsledder
- |
  bobsleigh
- |
  bobtail
- |
  bobtailed
- |
  bobwhite
- |
  Boccaccio
- |
  bocce
- |
  bocci
- |
  boccie
- |
  Bochum
- |
  bodacious
- |
  bodega
- |
  Bodhisattva
- |
  bodhisattva
- |
  bodice
- |
  bodied
- |
  bodiless
- |
  bodily
- |
  bodkin
- |
  bodyboard
- |
  bodyboarder
- |
  bodybuilder
- |
  bodybuilding
- |
  bodyguard
- |
  bodysuit
- |
  bodysurf
- |
  bodywork
- |
  Boeotia
- |
  Boeotian
- |
  Boethius
- |
  boffo
- |
  Bogart
- |
  bogey
- |
  bogeyman
- |
  boggle
- |
  boggy
- |
  bogie
- |
  Bogota
- |
  bogus
- |
  bogusly
- |
  bogusness
- |
  bogyman
- |
  Bohemia
- |
  Bohemian
- |
  bohemian
- |
  Bohemianism
- |
  bohemianism
- |
  Bohol
- |
  bohrium
- |
  boiler
- |
  boilermaker
- |
  boiling
- |
  Boise
- |
  boisterous
- |
  boisterously
- |
  bolas
- |
  boldface
- |
  boldfaced
- |
  boldly
- |
  boldness
- |
  bolero
- |
  Boleyn
- |
  Bolivar
- |
  bolivar
- |
  bolivares
- |
  Bolivia
- |
  Bolivian
- |
  boliviano
- |
  bollworm
- |
  Bologna
- |
  bologna
- |
  Bolognan
- |
  Bolognese
- |
  boloney
- |
  Bolshevik
- |
  Bolsheviki
- |
  Bolshevism
- |
  bolshevism
- |
  Bolshevist
- |
  Bolshoi
- |
  bolster
- |
  bolter
- |
  Bolton
- |
  bolus
- |
  bombard
- |
  bombardier
- |
  bombardment
- |
  bombast
- |
  bombastic
- |
  Bombay
- |
  bombazine
- |
  bombed
- |
  bomber
- |
  bombing
- |
  bombproof
- |
  bombshell
- |
  bombsight
- |
  bonanza
- |
  Bonaparte
- |
  bonbon
- |
  bondage
- |
  bondholder
- |
  bonding
- |
  bondman
- |
  bonds
- |
  bondservant
- |
  bondsman
- |
  bondswoman
- |
  bondwoman
- |
  boneblack
- |
  bonehead
- |
  boneless
- |
  boner
- |
  boney
- |
  bonfire
- |
  bongo
- |
  bongos
- |
  bonhomie
- |
  Boniface
- |
  boniness
- |
  Bonita
- |
  bonito
- |
  bonkers
- |
  bonnet
- |
  Bonnie
- |
  bonnie
- |
  bonny
- |
  bonobo
- |
  bonsai
- |
  bonus
- |
  bonze
- |
  booboo
- |
  booby
- |
  boodle
- |
  boogeyman
- |
  boogie
- |
  booing
- |
  bookbinder
- |
  bookbindery
- |
  bookbinding
- |
  bookcase
- |
  bookend
- |
  bookie
- |
  booking
- |
  bookish
- |
  bookkeeper
- |
  bookkeeping
- |
  booklet
- |
  bookmaker
- |
  bookmaking
- |
  bookmark
- |
  bookmarker
- |
  bookmobile
- |
  bookplate
- |
  books
- |
  bookseller
- |
  bookshelf
- |
  bookshelves
- |
  bookshop
- |
  bookstore
- |
  bookworm
- |
  Boolean
- |
  boombox
- |
  boomerang
- |
  booming
- |
  boondocks
- |
  boondoggle
- |
  boondoggler
- |
  Boone
- |
  boorish
- |
  boorishly
- |
  boorishness
- |
  boost
- |
  booster
- |
  boosterism
- |
  bootblack
- |
  bootee
- |
  Bootes
- |
  Booth
- |
  booth
- |
  Boothia
- |
  bootie
- |
  bootleg
- |
  bootlegger
- |
  bootlegging
- |
  bootless
- |
  bootlessly
- |
  bootlessness
- |
  bootlick
- |
  bootlicker
- |
  bootstrap
- |
  bootstraps
- |
  booty
- |
  booze
- |
  boozer
- |
  boozing
- |
  boozy
- |
  bopper
- |
  borate
- |
  borax
- |
  Bordeaux
- |
  bordello
- |
  Borden
- |
  border
- |
  borderland
- |
  borderline
- |
  Borders
- |
  Boreal
- |
  boreal
- |
  Boreas
- |
  bored
- |
  boredom
- |
  borer
- |
  Borges
- |
  Borgia
- |
  boring
- |
  boringly
- |
  Boris
- |
  borne
- |
  Bornean
- |
  Borneo
- |
  Borodin
- |
  boron
- |
  borough
- |
  borrow
- |
  borrower
- |
  borrowing
- |
  borrowings
- |
  borsch
- |
  borscht
- |
  borsht
- |
  borzoi
- |
  boscage
- |
  Bosch
- |
  boskage
- |
  bosky
- |
  Bosnia
- |
  Bosnian
- |
  bosom
- |
  bosomed
- |
  bosomy
- |
  boson
- |
  Bosporus
- |
  bossiness
- |
  bossism
- |
  bossy
- |
  Boston
- |
  Bostonian
- |
  bosun
- |
  Boswell
- |
  botanic
- |
  botanical
- |
  botanicals
- |
  botanist
- |
  botanize
- |
  botany
- |
  botch
- |
  botcher
- |
  botchily
- |
  botchy
- |
  botfly
- |
  bother
- |
  bothered
- |
  bothersome
- |
  Bothnia
- |
  Botswana
- |
  Botticelli
- |
  bottle
- |
  bottled
- |
  bottleful
- |
  bottleneck
- |
  bottler
- |
  bottom
- |
  bottomland
- |
  bottomless
- |
  bottoms
- |
  botulism
- |
  Boudicca
- |
  boudoir
- |
  bouffant
- |
  bough
- |
  bought
- |
  bouillon
- |
  Boulder
- |
  boulder
- |
  bouldered
- |
  boulevard
- |
  Boulez
- |
  bounce
- |
  bouncer
- |
  bouncily
- |
  bouncing
- |
  bouncy
- |
  bound
- |
  boundary
- |
  bounden
- |
  bounder
- |
  boundless
- |
  boundlessly
- |
  bounds
- |
  bounteous
- |
  bounteously
- |
  bountiful
- |
  bountifully
- |
  bounty
- |
  bouquet
- |
  Bourbon
- |
  bourbon
- |
  bourgeois
- |
  bourgeoisie
- |
  bourgeoisify
- |
  Bourgogne
- |
  bourn
- |
  bourne
- |
  Bournemouth
- |
  Bourse
- |
  bourse
- |
  boutique
- |
  boutonniere
- |
  bovine
- |
  bovinely
- |
  bowdlerism
- |
  bowdlerize
- |
  bowdlerized
- |
  bowel
- |
  bowels
- |
  bower
- |
  Bowery
- |
  Bowie
- |
  bowknot
- |
  bowlder
- |
  bowleg
- |
  bowlegged
- |
  bowlegs
- |
  bowler
- |
  bowlful
- |
  bowline
- |
  bowling
- |
  bowllike
- |
  bowls
- |
  bowman
- |
  bowsprit
- |
  bowstring
- |
  boxcar
- |
  boxer
- |
  boxful
- |
  boxing
- |
  boxlike
- |
  boxwood
- |
  boycott
- |
  boyfriend
- |
  boyhood
- |
  boyish
- |
  boyishly
- |
  boyishness
- |
  Boyle
- |
  boysenberry
- |
  brace
- |
  bracelet
- |
  bracero
- |
  braces
- |
  brachial
- |
  brachiate
- |
  brachiation
- |
  brachiator
- |
  brachiosaur
- |
  bracing
- |
  bracken
- |
  bracket
- |
  brackish
- |
  brackishness
- |
  bract
- |
  Bradbury
- |
  Braddock
- |
  Bradford
- |
  Bradley
- |
  Bradstreet
- |
  Brady
- |
  braggadocio
- |
  braggart
- |
  bragger
- |
  Brahe
- |
  Brahma
- |
  Brahman
- |
  Brahmanic
- |
  Brahmanical
- |
  Brahmanism
- |
  Brahmanist
- |
  Brahmaputra
- |
  Brahmin
- |
  Brahminic
- |
  Brahminical
- |
  Brahminism
- |
  Brahms
- |
  Brahmsian
- |
  braid
- |
  braided
- |
  braider
- |
  braiding
- |
  Braila
- |
  Braille
- |
  braille
- |
  brain
- |
  brainchild
- |
  brained
- |
  braininess
- |
  brainless
- |
  brainpower
- |
  brains
- |
  brainstorm
- |
  brainteaser
- |
  brainwash
- |
  brainwashing
- |
  brainy
- |
  braise
- |
  brake
- |
  brakeless
- |
  brakeman
- |
  braless
- |
  bramble
- |
  brambly
- |
  Brampton
- |
  branch
- |
  branched
- |
  branchless
- |
  branchlike
- |
  brand
- |
  Brandeis
- |
  Brandenburg
- |
  brander
- |
  brandish
- |
  brandisher
- |
  brandless
- |
  Brando
- |
  Brandon
- |
  Brandt
- |
  Brandy
- |
  brandy
- |
  Brant
- |
  brant
- |
  Braque
- |
  brash
- |
  brashly
- |
  brashness
- |
  Brasilia
- |
  Brasov
- |
  brass
- |
  brasserie
- |
  brasses
- |
  brassiere
- |
  brassily
- |
  brassiness
- |
  brassy
- |
  Bratislava
- |
  brattiness
- |
  bratty
- |
  bratwurst
- |
  Braun
- |
  bravado
- |
  brave
- |
  bravely
- |
  braveness
- |
  bravery
- |
  bravo
- |
  bravura
- |
  brawl
- |
  brawler
- |
  brawling
- |
  brawn
- |
  brawniness
- |
  brawny
- |
  braze
- |
  brazen
- |
  brazenly
- |
  brazenness
- |
  brazer
- |
  brazier
- |
  Brazil
- |
  Brazilian
- |
  Brazos
- |
  Brazzaville
- |
  breach
- |
  bread
- |
  breadbasket
- |
  breadboard
- |
  breadcrumb
- |
  breadcrumbs
- |
  breaded
- |
  breadfruit
- |
  breadstuff
- |
  breadth
- |
  breadwinner
- |
  break
- |
  breakable
- |
  breakage
- |
  breakaway
- |
  breakdown
- |
  breaker
- |
  breakfast
- |
  breakfront
- |
  breakneck
- |
  breakout
- |
  breakthrough
- |
  breakup
- |
  breakwater
- |
  bream
- |
  breast
- |
  breastbone
- |
  breastplate
- |
  breaststroke
- |
  breastwork
- |
  breath
- |
  breathable
- |
  breathalyze
- |
  Breathalyzer
- |
  breathe
- |
  breather
- |
  breathing
- |
  breathless
- |
  breathlessly
- |
  breathtaking
- |
  breathy
- |
  breccia
- |
  Brecht
- |
  Brechtian
- |
  Breda
- |
  breech
- |
  breechcloth
- |
  breeches
- |
  breed
- |
  breeder
- |
  breeding
- |
  breeze
- |
  breezeless
- |
  breezeway
- |
  breezily
- |
  breeziness
- |
  breezy
- |
  Bremen
- |
  Bremerhaven
- |
  Brenda
- |
  Brendan
- |
  Brenner
- |
  Brent
- |
  Brescia
- |
  Brest
- |
  Brethren
- |
  brethren
- |
  Breton
- |
  Brett
- |
  Breughel
- |
  breve
- |
  brevet
- |
  breviary
- |
  brevity
- |
  brewer
- |
  brewery
- |
  brewing
- |
  brewpub
- |
  Breyer
- |
  Brezhnev
- |
  Brian
- |
  briar
- |
  bribable
- |
  bribe
- |
  briber
- |
  bribery
- |
  Brice
- |
  brick
- |
  brickbat
- |
  bricklayer
- |
  bricklaying
- |
  bricolage
- |
  bridal
- |
  Bridalveil
- |
  bride
- |
  bridegroom
- |
  bridesmaid
- |
  bridge
- |
  bridgeable
- |
  bridgehead
- |
  Bridgeport
- |
  Bridger
- |
  Bridges
- |
  Bridget
- |
  Bridgetown
- |
  bridgework
- |
  bridle
- |
  brief
- |
  briefcase
- |
  briefing
- |
  briefly
- |
  briefness
- |
  briefs
- |
  brier
- |
  briery
- |
  brigade
- |
  brigadier
- |
  brigand
- |
  brigandage
- |
  brigandry
- |
  brigantine
- |
  bright
- |
  brighten
- |
  brightener
- |
  brightly
- |
  brightness
- |
  Brighton
- |
  brights
- |
  Brigitte
- |
  brill
- |
  brilliance
- |
  brilliancy
- |
  brilliant
- |
  brilliantine
- |
  brilliantly
- |
  brimful
- |
  brimless
- |
  brimstone
- |
  brindle
- |
  brindled
- |
  brine
- |
  bring
- |
  bringer
- |
  brininess
- |
  brink
- |
  brinkmanship
- |
  briny
- |
  brioche
- |
  briquet
- |
  briquette
- |
  Brisbane
- |
  brisk
- |
  brisket
- |
  briskly
- |
  briskness
- |
  brisling
- |
  bristle
- |
  bristlelike
- |
  bristly
- |
  Bristol
- |
  Britain
- |
  Britannia
- |
  Britannic
- |
  britches
- |
  Briticism
- |
  British
- |
  Britishism
- |
  Britishness
- |
  Briton
- |
  Brittany
- |
  Britten
- |
  brittle
- |
  brittlely
- |
  brittleness
- |
  broach
- |
  broacher
- |
  broad
- |
  broadband
- |
  broadcast
- |
  broadcaster
- |
  broadcasting
- |
  broadcloth
- |
  broaden
- |
  broadener
- |
  broadloom
- |
  broadly
- |
  broadminded
- |
  broadness
- |
  broadsheet
- |
  broadside
- |
  broadsword
- |
  broadtail
- |
  Broadway
- |
  brocade
- |
  broccoli
- |
  brochette
- |
  brochure
- |
  Brockton
- |
  Brodsky
- |
  brogan
- |
  brogue
- |
  broil
- |
  broiler
- |
  broiling
- |
  broke
- |
  broken
- |
  brokenly
- |
  brokenness
- |
  broker
- |
  brokerage
- |
  broking
- |
  bromeliad
- |
  bromide
- |
  bromidic
- |
  bromine
- |
  Bromley
- |
  bronc
- |
  bronchi
- |
  bronchial
- |
  bronchitic
- |
  bronchitis
- |
  broncho
- |
  bronchus
- |
  bronco
- |
  broncobuster
- |
  Bronte
- |
  brontosaur
- |
  brontosaurus
- |
  Bronx
- |
  bronze
- |
  bronzy
- |
  brooch
- |
  brood
- |
  brooder
- |
  brooding
- |
  broodingly
- |
  broodmare
- |
  broody
- |
  brook
- |
  Brooke
- |
  brooklet
- |
  Brooklyn
- |
  Brooks
- |
  broom
- |
  broomstick
- |
  broth
- |
  brothel
- |
  brother
- |
  brotherhood
- |
  brotherly
- |
  brougham
- |
  brought
- |
  brouhaha
- |
  browbeat
- |
  browbeaten
- |
  Brown
- |
  brown
- |
  Browne
- |
  brownfield
- |
  Brownie
- |
  brownie
- |
  Brownies
- |
  Browning
- |
  brownish
- |
  brownness
- |
  brownout
- |
  brownstone
- |
  Brownsville
- |
  browse
- |
  browser
- |
  Bruce
- |
  Bruckner
- |
  Bruegel
- |
  Brueghel
- |
  Bruges
- |
  Brugge
- |
  bruin
- |
  bruise
- |
  bruised
- |
  bruiser
- |
  bruising
- |
  bruit
- |
  brunch
- |
  Brunei
- |
  Bruneian
- |
  Brunelleschi
- |
  brunet
- |
  brunette
- |
  Brunnhilde
- |
  Bruno
- |
  Brunswick
- |
  brunt
- |
  brush
- |
  brushoff
- |
  brushwood
- |
  brushwork
- |
  brushy
- |
  brusk
- |
  brusque
- |
  brusquely
- |
  brusqueness
- |
  brusquerie
- |
  Brussels
- |
  brutal
- |
  brutalism
- |
  brutalist
- |
  brutality
- |
  brutalize
- |
  brutally
- |
  brute
- |
  brutish
- |
  brutishly
- |
  brutishness
- |
  Brutus
- |
  Bryan
- |
  Bryansk
- |
  Bryant
- |
  Bryce
- |
  Brynner
- |
  bubba
- |
  bubble
- |
  bubblegum
- |
  bubbly
- |
  Buber
- |
  Bucaramanga
- |
  buccal
- |
  buccaneer
- |
  buccaneering
- |
  Buchanan
- |
  Bucharest
- |
  buckboard
- |
  bucker
- |
  bucket
- |
  bucketful
- |
  buckeye
- |
  Buckingham
- |
  buckle
- |
  buckler
- |
  buckram
- |
  bucksaw
- |
  buckshot
- |
  buckskin
- |
  buckskins
- |
  buckteeth
- |
  bucktooth
- |
  bucktoothed
- |
  buckwheat
- |
  buckyball
- |
  bucolic
- |
  bucolically
- |
  Budapest
- |
  budder
- |
  Buddha
- |
  Buddhism
- |
  Buddhist
- |
  budding
- |
  Buddy
- |
  buddy
- |
  budge
- |
  budgerigar
- |
  budget
- |
  budgetary
- |
  budgeting
- |
  budgie
- |
  budlike
- |
  Buffalo
- |
  buffalo
- |
  buffer
- |
  buffered
- |
  buffet
- |
  buffeter
- |
  buffeting
- |
  buffing
- |
  Buffon
- |
  buffoon
- |
  buffoonery
- |
  buffoonish
- |
  Buford
- |
  bugaboo
- |
  bugbear
- |
  bugger
- |
  buggery
- |
  bugging
- |
  buggy
- |
  bugle
- |
  bugler
- |
  build
- |
  builder
- |
  building
- |
  buildup
- |
  built
- |
  Bujumbura
- |
  Bukharin
- |
  Bukovina
- |
  Bulawayo
- |
  bulbous
- |
  Bulfinch
- |
  Bulganin
- |
  Bulgar
- |
  Bulgaria
- |
  Bulgarian
- |
  bulge
- |
  bulghur
- |
  bulginess
- |
  bulgur
- |
  bulgy
- |
  bulimarexia
- |
  bulimarexic
- |
  bulimia
- |
  bulimic
- |
  bulkhead
- |
  bulkily
- |
  bulkiness
- |
  bulky
- |
  bulldog
- |
  bulldoze
- |
  bulldozer
- |
  bullet
- |
  bulletin
- |
  bulletproof
- |
  bullfight
- |
  bullfighter
- |
  bullfighting
- |
  bullfinch
- |
  bullfrog
- |
  bullhead
- |
  bullheaded
- |
  bullheadedly
- |
  bullhorn
- |
  bullion
- |
  bullish
- |
  bullishly
- |
  bullishness
- |
  bullock
- |
  bullpen
- |
  bullring
- |
  bullshit
- |
  bullshitter
- |
  bullwhip
- |
  bully
- |
  bullying
- |
  bullyrag
- |
  bulrush
- |
  Bultmann
- |
  bulwark
- |
  bulwarks
- |
  bumble
- |
  bumblebee
- |
  bumbler
- |
  bumbling
- |
  bummed
- |
  bummer
- |
  bumper
- |
  bumpiness
- |
  bumpkin
- |
  Bumppo
- |
  bumptious
- |
  bumptiously
- |
  bumpy
- |
  bunch
- |
  Bunche
- |
  bunchy
- |
  bunco
- |
  buncombe
- |
  Bundestag
- |
  bundle
- |
  bundling
- |
  Bundt
- |
  bungalow
- |
  bungee
- |
  bunghole
- |
  bungle
- |
  bungler
- |
  bungling
- |
  Bunin
- |
  bunion
- |
  Bunker
- |
  bunker
- |
  bunkhouse
- |
  bunko
- |
  bunkum
- |
  bunny
- |
  bunter
- |
  bunting
- |
  Bunuel
- |
  Bunyan
- |
  buoyancy
- |
  buoyant
- |
  buoyantly
- |
  Burbank
- |
  burbs
- |
  burden
- |
  burdened
- |
  burdensome
- |
  burdock
- |
  bureau
- |
  bureaucracy
- |
  bureaucrat
- |
  bureaucratic
- |
  bureaux
- |
  buret
- |
  burette
- |
  burgeon
- |
  burgeoning
- |
  burger
- |
  Burgess
- |
  burgess
- |
  burgh
- |
  burghal
- |
  burgher
- |
  burglar
- |
  burglarize
- |
  burglarproof
- |
  burglary
- |
  burgle
- |
  burgomaster
- |
  Burgos
- |
  Burgoyne
- |
  Burgundian
- |
  Burgundy
- |
  burgundy
- |
  burial
- |
  Burke
- |
  burlap
- |
  burled
- |
  burlesque
- |
  burley
- |
  burliness
- |
  Burlington
- |
  burly
- |
  Burma
- |
  Burman
- |
  Burmese
- |
  burnable
- |
  Burnaby
- |
  burner
- |
  Burnett
- |
  burning
- |
  burnish
- |
  burnished
- |
  burnisher
- |
  burnishing
- |
  burnoose
- |
  burnous
- |
  burnout
- |
  Burns
- |
  Burnsian
- |
  Burnside
- |
  burnt
- |
  burrito
- |
  burro
- |
  Burroughs
- |
  burrow
- |
  burrower
- |
  burry
- |
  Bursa
- |
  bursa
- |
  bursae
- |
  bursar
- |
  bursary
- |
  bursitis
- |
  burst
- |
  bursting
- |
  Burton
- |
  Burundi
- |
  Burundian
- |
  busboy
- |
  busby
- |
  busgirl
- |
  bushed
- |
  bushel
- |
  bushido
- |
  bushily
- |
  bushiness
- |
  bushing
- |
  Bushman
- |
  bushman
- |
  bushmaster
- |
  bushwhack
- |
  bushwhacker
- |
  bushy
- |
  busily
- |
  business
- |
  businesslike
- |
  businessman
- |
  busing
- |
  busker
- |
  buskin
- |
  buskined
- |
  busman
- |
  busses
- |
  bussing
- |
  busted
- |
  buster
- |
  bustle
- |
  bustler
- |
  busybody
- |
  busyness
- |
  busywork
- |
  butadiene
- |
  butane
- |
  butch
- |
  butcher
- |
  butcherer
- |
  butchery
- |
  buteo
- |
  Butler
- |
  butler
- |
  Butte
- |
  butte
- |
  butter
- |
  buttercup
- |
  butterfat
- |
  butterfish
- |
  butterflies
- |
  butterfly
- |
  buttermilk
- |
  butternut
- |
  butterscotch
- |
  buttery
- |
  buttock
- |
  buttocks
- |
  button
- |
  buttonhole
- |
  buttress
- |
  buttressed
- |
  butut
- |
  butyl
- |
  buxom
- |
  buxomness
- |
  buyback
- |
  buyer
- |
  buyout
- |
  buzzard
- |
  buzzer
- |
  buzzing
- |
  buzzsaw
- |
  buzzword
- |
  Bydgoszcz
- |
  Byelarus
- |
  byelaw
- |
  Byelorussia
- |
  Byelorussian
- |
  bygone
- |
  bygones
- |
  bylaw
- |
  byline
- |
  byliner
- |
  bypass
- |
  bypath
- |
  byplay
- |
  byproduct
- |
  byroad
- |
  Byron
- |
  Byronic
- |
  bystander
- |
  byway
- |
  byword
- |
  Byzantine
- |
  byzantine
- |
  Byzantinism
- |
  Byzantium
- |
  cabal
- |
  Cabala
- |
  cabala
- |
  caballero
- |
  cabana
- |
  cabaret
- |
  cabbage
- |
  cabbagy
- |
  Cabbala
- |
  cabbie
- |
  cabby
- |
  cabernet
- |
  cabin
- |
  Cabinet
- |
  cabinet
- |
  cabinetmaker
- |
  cabinetry
- |
  cabinetwork
- |
  cable
- |
  cablecast
- |
  cablegram
- |
  cablevision
- |
  cabochon
- |
  caboodle
- |
  caboose
- |
  Cabot
- |
  cabotage
- |
  Cabrini
- |
  cabriolet
- |
  cabstand
- |
  cacao
- |
  cacciatore
- |
  cachalot
- |
  cache
- |
  cachepot
- |
  cachet
- |
  cachexia
- |
  cachinnate
- |
  cachinnation
- |
  cacique
- |
  cackle
- |
  cackler
- |
  cacodemon
- |
  cacoethes
- |
  cacophonous
- |
  cacophony
- |
  cacti
- |
  cactus
- |
  cadastral
- |
  cadaver
- |
  cadaverous
- |
  cadaverously
- |
  caddie
- |
  caddish
- |
  caddishly
- |
  caddishness
- |
  Caddoan
- |
  caddy
- |
  cadence
- |
  cadenced
- |
  cadency
- |
  cadenza
- |
  cadet
- |
  cadetship
- |
  Cadette
- |
  cadge
- |
  cadger
- |
  Cadillac
- |
  Cadiz
- |
  cadmic
- |
  cadmium
- |
  cadre
- |
  caducei
- |
  caduceus
- |
  caducity
- |
  caeca
- |
  caecum
- |
  Caedmon
- |
  Caelum
- |
  Caernarvon
- |
  Caesar
- |
  caesar
- |
  Caesarea
- |
  Caesarean
- |
  caesarean
- |
  Caesarian
- |
  caesarian
- |
  caesium
- |
  caesura
- |
  caesurae
- |
  caesural
- |
  cafeteria
- |
  caffein
- |
  caffeinated
- |
  caffeine
- |
  caftan
- |
  cager
- |
  cagey
- |
  cagily
- |
  caginess
- |
  Cagliari
- |
  Cagney
- |
  Caguas
- |
  cahoot
- |
  cahoots
- |
  caiman
- |
  Caine
- |
  Cainozoic
- |
  Cairene
- |
  cairn
- |
  Cairo
- |
  caisson
- |
  caitiff
- |
  Caitlin
- |
  Cajan
- |
  cajole
- |
  cajolement
- |
  cajoler
- |
  cajolery
- |
  cajolingly
- |
  Cajun
- |
  cakewalk
- |
  cakey
- |
  calabash
- |
  calaboose
- |
  Calabria
- |
  Calabrian
- |
  caladium
- |
  Calais
- |
  calamari
- |
  calamine
- |
  calamitous
- |
  calamitously
- |
  calamity
- |
  calcareous
- |
  calces
- |
  calciferous
- |
  calcific
- |
  calcify
- |
  calcimine
- |
  calcination
- |
  calcine
- |
  calcite
- |
  calcitic
- |
  calcium
- |
  calculable
- |
  calculate
- |
  calculated
- |
  calculatedly
- |
  calculating
- |
  calculation
- |
  calculative
- |
  calculator
- |
  calculi
- |
  calculus
- |
  Calcutta
- |
  Calcuttan
- |
  Calder
- |
  caldera
- |
  caldron
- |
  Caleb
- |
  Caledonia
- |
  Caledonian
- |
  calendar
- |
  calender
- |
  calendric
- |
  calendrical
- |
  calends
- |
  calendula
- |
  calfskin
- |
  Calgary
- |
  Calhoun
- |
  caliber
- |
  calibrate
- |
  calibration
- |
  calibrator
- |
  calibre
- |
  calices
- |
  calico
- |
  calif
- |
  California
- |
  Californian
- |
  californium
- |
  Caligula
- |
  caliper
- |
  calipers
- |
  caliph
- |
  caliphate
- |
  calisthenic
- |
  calisthenics
- |
  calix
- |
  calker
- |
  calla
- |
  Callaghan
- |
  Callao
- |
  Callas
- |
  callback
- |
  called
- |
  caller
- |
  calligrapher
- |
  calligraphic
- |
  calligraphy
- |
  calling
- |
  Calliope
- |
  calliope
- |
  calliper
- |
  callipers
- |
  callipygean
- |
  callipygian
- |
  callipygous
- |
  callosity
- |
  callous
- |
  calloused
- |
  callously
- |
  callousness
- |
  callow
- |
  callowly
- |
  callowness
- |
  callus
- |
  callused
- |
  calmative
- |
  calming
- |
  calmly
- |
  calmness
- |
  calomel
- |
  Caloocan
- |
  caloric
- |
  calorically
- |
  calorie
- |
  calorific
- |
  calorimeter
- |
  calorimetry
- |
  calque
- |
  calumet
- |
  calumniate
- |
  calumniation
- |
  calumniator
- |
  calumnious
- |
  calumniously
- |
  calumny
- |
  calvados
- |
  Calvary
- |
  calvary
- |
  calve
- |
  Calvert
- |
  calves
- |
  Calvin
- |
  Calvinism
- |
  Calvinist
- |
  Calvinistic
- |
  calvities
- |
  calyces
- |
  Calypso
- |
  calypso
- |
  Calypsonian
- |
  calyx
- |
  calzone
- |
  Camaguey
- |
  camaraderie
- |
  camber
- |
  cambia
- |
  cambial
- |
  cambium
- |
  Cambodia
- |
  Cambodian
- |
  Cambria
- |
  Cambrian
- |
  cambric
- |
  Cambridge
- |
  camcorder
- |
  Camden
- |
  camel
- |
  camelhair
- |
  camellia
- |
  Camelot
- |
  Camembert
- |
  cameo
- |
  camera
- |
  cameraman
- |
  camerawoman
- |
  Cameron
- |
  Cameroon
- |
  Cameroonian
- |
  Cameroun
- |
  Camiguin
- |
  Camilla
- |
  Camille
- |
  camisole
- |
  Camoens
- |
  Camoes
- |
  camomile
- |
  camouflage
- |
  camouflager
- |
  campaign
- |
  campaigner
- |
  Campania
- |
  campanile
- |
  campanili
- |
  campanology
- |
  Campeche
- |
  camped
- |
  camper
- |
  campesino
- |
  Campfire
- |
  campfire
- |
  campground
- |
  camphor
- |
  camphorated
- |
  campily
- |
  Campinas
- |
  campiness
- |
  camping
- |
  Campion
- |
  camporee
- |
  Campos
- |
  campsite
- |
  campus
- |
  campy
- |
  camshaft
- |
  Camus
- |
  Canaan
- |
  Canaanite
- |
  Canada
- |
  Canadian
- |
  Canadianism
- |
  canaille
- |
  canal
- |
  Canaletto
- |
  canalization
- |
  canalize
- |
  canape
- |
  canard
- |
  Canary
- |
  canary
- |
  canasta
- |
  Canaveral
- |
  Canberra
- |
  cancan
- |
  cancel
- |
  cancelable
- |
  canceler
- |
  cancellation
- |
  canceller
- |
  Cancer
- |
  cancer
- |
  cancerous
- |
  cancerously
- |
  Cancun
- |
  Candace
- |
  candela
- |
  candelabra
- |
  candelabrum
- |
  candescence
- |
  candescent
- |
  Candia
- |
  candid
- |
  candidacy
- |
  candidate
- |
  candidature
- |
  Candide
- |
  candidly
- |
  candidness
- |
  candied
- |
  candle
- |
  candlelight
- |
  candlelit
- |
  Candlemas
- |
  candlepin
- |
  candlepower
- |
  candler
- |
  candlestick
- |
  candlewick
- |
  candor
- |
  candour
- |
  candy
- |
  candystriper
- |
  candytuft
- |
  canebrake
- |
  caner
- |
  canine
- |
  canister
- |
  canker
- |
  cankerous
- |
  cankerworm
- |
  canna
- |
  cannabis
- |
  canned
- |
  cannelloni
- |
  canner
- |
  cannery
- |
  Cannes
- |
  cannibal
- |
  cannibalism
- |
  cannibalize
- |
  cannily
- |
  canniness
- |
  Canning
- |
  cannoli
- |
  cannon
- |
  cannonade
- |
  cannonball
- |
  cannoneer
- |
  cannonfodder
- |
  cannot
- |
  cannula
- |
  cannulae
- |
  canny
- |
  canoe
- |
  canoeist
- |
  canola
- |
  canon
- |
  canonic
- |
  canonical
- |
  canonically
- |
  canonicity
- |
  canonization
- |
  canonize
- |
  canopied
- |
  Canopus
- |
  canopy
- |
  Canova
- |
  canst
- |
  cantabile
- |
  cantaloup
- |
  cantaloupe
- |
  cantankerous
- |
  cantata
- |
  canteen
- |
  canteloupe
- |
  canter
- |
  Canterbury
- |
  canthi
- |
  canthus
- |
  canticle
- |
  Canticles
- |
  cantilever
- |
  cantilevered
- |
  cantina
- |
  cantingly
- |
  cantle
- |
  canto
- |
  Canton
- |
  canton
- |
  cantonal
- |
  Cantonese
- |
  cantonment
- |
  cantor
- |
  cantorial
- |
  Canute
- |
  canvas
- |
  canvasback
- |
  canvass
- |
  canvasser
- |
  canyon
- |
  caoutchouc
- |
  capability
- |
  capable
- |
  capably
- |
  capacious
- |
  capaciously
- |
  capacitance
- |
  capacitate
- |
  capacitative
- |
  capacitive
- |
  capacitor
- |
  capacity
- |
  caparison
- |
  caped
- |
  Capella
- |
  caper
- |
  capeskin
- |
  Capet
- |
  Capetown
- |
  capful
- |
  capillarity
- |
  capillary
- |
  capital
- |
  capitalise
- |
  capitalism
- |
  capitalist
- |
  capitalistic
- |
  capitalize
- |
  capitally
- |
  capitation
- |
  Capitol
- |
  capitol
- |
  capitulate
- |
  capitulation
- |
  capitulator
- |
  capitulatory
- |
  caplet
- |
  capon
- |
  Capone
- |
  Capote
- |
  Cappadocia
- |
  Cappadocian
- |
  capping
- |
  cappuccino
- |
  Capra
- |
  Capri
- |
  capriccio
- |
  caprice
- |
  capricious
- |
  capriciously
- |
  Capricorn
- |
  Capricornis
- |
  capriole
- |
  capsful
- |
  capsicum
- |
  capsid
- |
  capsize
- |
  capstan
- |
  capstone
- |
  capsular
- |
  capsulate
- |
  capsulated
- |
  capsulation
- |
  capsule
- |
  capsulize
- |
  Captain
- |
  captain
- |
  captaincy
- |
  captainship
- |
  caption
- |
  captious
- |
  captiously
- |
  captiousness
- |
  captivate
- |
  captivating
- |
  captivation
- |
  captivator
- |
  captive
- |
  captivity
- |
  captor
- |
  capture
- |
  Capuchin
- |
  capuchin
- |
  capybara
- |
  carabiner
- |
  Caracalla
- |
  Caracas
- |
  caracole
- |
  caracul
- |
  carafe
- |
  carambola
- |
  caramel
- |
  caramelize
- |
  carapace
- |
  carat
- |
  Caravaggio
- |
  caravan
- |
  caravansary
- |
  caravanserai
- |
  caravansery
- |
  caravel
- |
  caravelle
- |
  caraway
- |
  carbide
- |
  carbine
- |
  carbohydrate
- |
  carbolic
- |
  carbon
- |
  carbonaceous
- |
  carbonate
- |
  carbonated
- |
  carbonation
- |
  carbonic
- |
  carbonize
- |
  carbonous
- |
  Carborundum
- |
  carborundum
- |
  carboy
- |
  carbuncle
- |
  carbuncular
- |
  carburet
- |
  carburetion
- |
  carburetor
- |
  carburetter
- |
  carburettor
- |
  carburize
- |
  carcase
- |
  carcass
- |
  carcinogen
- |
  carcinogenic
- |
  carcinoma
- |
  carcinomata
- |
  cardamom
- |
  cardamon
- |
  cardboard
- |
  carder
- |
  cardiac
- |
  Cardiff
- |
  cardigan
- |
  cardinal
- |
  cardinalate
- |
  cardinally
- |
  cardinalship
- |
  cardiogram
- |
  cardiograph
- |
  cardiography
- |
  cardiologist
- |
  cardiology
- |
  cards
- |
  cardsharp
- |
  cardsharper
- |
  cardsharping
- |
  careen
- |
  careener
- |
  career
- |
  careerism
- |
  careerist
- |
  carefree
- |
  careful
- |
  carefully
- |
  carefulness
- |
  caregiver
- |
  caregiving
- |
  careless
- |
  carelessly
- |
  carelessness
- |
  carer
- |
  caress
- |
  caresser
- |
  caret
- |
  caretaker
- |
  careworn
- |
  Carey
- |
  carfare
- |
  cargo
- |
  carhop
- |
  Carib
- |
  Cariban
- |
  Caribbean
- |
  caribou
- |
  caricatural
- |
  caricature
- |
  caricaturist
- |
  caries
- |
  carillon
- |
  Carina
- |
  caring
- |
  carious
- |
  caritas
- |
  carjack
- |
  carjacker
- |
  carjacking
- |
  Carla
- |
  Carlene
- |
  Carleton
- |
  Carlisle
- |
  carload
- |
  Carlos
- |
  Carlotta
- |
  Carlyle
- |
  Carmarthen
- |
  Carmel
- |
  Carmen
- |
  Carmichael
- |
  carminative
- |
  Carmine
- |
  carmine
- |
  carnage
- |
  carnal
- |
  carnality
- |
  carnally
- |
  carnation
- |
  carnauba
- |
  Carne
- |
  Carnegie
- |
  carnelian
- |
  carney
- |
  carnie
- |
  carnival
- |
  carnivora
- |
  carnivore
- |
  carnivorous
- |
  carny
- |
  carob
- |
  Carol
- |
  carol
- |
  Carole
- |
  caroler
- |
  Carolina
- |
  Carolinas
- |
  Caroline
- |
  Carolinian
- |
  caroller
- |
  Carolyn
- |
  carom
- |
  carotene
- |
  carotid
- |
  carousal
- |
  carouse
- |
  carousel
- |
  carouser
- |
  carousing
- |
  carpal
- |
  carpark
- |
  Carpathian
- |
  carpel
- |
  carpenter
- |
  carpentry
- |
  carper
- |
  carpet
- |
  carpetbag
- |
  carpetbagger
- |
  carpeting
- |
  carpi
- |
  carping
- |
  carpool
- |
  carpooling
- |
  carport
- |
  carpus
- |
  Carracci
- |
  carrageen
- |
  carrageenan
- |
  carrageenin
- |
  carragheen
- |
  carrel
- |
  carrell
- |
  Carreras
- |
  carriage
- |
  carriageway
- |
  Carrie
- |
  carrier
- |
  carrion
- |
  Carroll
- |
  carrot
- |
  carrousel
- |
  carry
- |
  carryall
- |
  carryon
- |
  carryout
- |
  carryover
- |
  carsick
- |
  carsickness
- |
  Carson
- |
  cartage
- |
  Cartagena
- |
  cartel
- |
  cartelism
- |
  Carter
- |
  carter
- |
  Cartesian
- |
  Cartesianism
- |
  Carthage
- |
  Carthaginian
- |
  Cartier
- |
  cartilage
- |
  cartographer
- |
  cartographic
- |
  cartography
- |
  cartomancy
- |
  carton
- |
  cartoon
- |
  cartoonish
- |
  cartoonist
- |
  cartoony
- |
  cartouche
- |
  cartridge
- |
  cartwheel
- |
  Cartwright
- |
  caruncle
- |
  caruncular
- |
  Caruso
- |
  carve
- |
  carvel
- |
  Carver
- |
  carver
- |
  carving
- |
  carwash
- |
  caryatid
- |
  caryatides
- |
  Caryl
- |
  casaba
- |
  Casablanca
- |
  Casals
- |
  Casanova
- |
  cascade
- |
  Cascades
- |
  cascara
- |
  caseharden
- |
  casein
- |
  caseload
- |
  casemate
- |
  casement
- |
  casette
- |
  casework
- |
  caseworker
- |
  cashbook
- |
  cashew
- |
  cashflow
- |
  cashier
- |
  cashiered
- |
  Cashmere
- |
  cashmere
- |
  casing
- |
  casino
- |
  casket
- |
  Casper
- |
  casque
- |
  Cassandra
- |
  Cassatt
- |
  cassava
- |
  casserole
- |
  cassette
- |
  cassia
- |
  cassino
- |
  Cassiopeia
- |
  cassiterite
- |
  Cassius
- |
  cassock
- |
  cassowary
- |
  castanet
- |
  castanets
- |
  castaway
- |
  caste
- |
  castellated
- |
  caster
- |
  castigate
- |
  castigation
- |
  castigator
- |
  castigatory
- |
  Castile
- |
  Castilian
- |
  Castilla
- |
  casting
- |
  castle
- |
  Castlereagh
- |
  castoff
- |
  Castor
- |
  castor
- |
  castrate
- |
  castrater
- |
  castration
- |
  castrator
- |
  Castries
- |
  Castro
- |
  casual
- |
  casually
- |
  casualness
- |
  casualty
- |
  casuist
- |
  casuistic
- |
  casuistical
- |
  casuistry
- |
  catabolic
- |
  catabolism
- |
  catachreses
- |
  catachresis
- |
  catachrestic
- |
  cataclysm
- |
  cataclysmal
- |
  cataclysmic
- |
  catacomb
- |
  catacombs
- |
  catafalque
- |
  Catalan
- |
  catalepsy
- |
  cataleptic
- |
  catalog
- |
  cataloger
- |
  catalogue
- |
  cataloguer
- |
  Catalonia
- |
  Catalonian
- |
  catalpa
- |
  catalyses
- |
  catalysis
- |
  catalyst
- |
  catalytic
- |
  catalyze
- |
  catalyzer
- |
  catamaran
- |
  catamite
- |
  catamount
- |
  Catanduanes
- |
  Catania
- |
  catapult
- |
  cataract
- |
  catarrh
- |
  catarrhal
- |
  catastrophe
- |
  catastrophic
- |
  catatonia
- |
  catatonic
- |
  Catawba
- |
  catbird
- |
  catboat
- |
  catcall
- |
  catch
- |
  catchall
- |
  catcher
- |
  catchiness
- |
  catching
- |
  catchment
- |
  catchpenny
- |
  catchup
- |
  catchword
- |
  catchy
- |
  catechetic
- |
  catechetical
- |
  catechetics
- |
  catechise
- |
  catechism
- |
  catechismal
- |
  catechist
- |
  catechize
- |
  catechizer
- |
  catechumen
- |
  categoric
- |
  categorical
- |
  categorise
- |
  categorize
- |
  category
- |
  catenary
- |
  catenated
- |
  catenation
- |
  cater
- |
  catercorner
- |
  caterer
- |
  catering
- |
  caterpillar
- |
  caterwaul
- |
  caterwauling
- |
  catfish
- |
  catgut
- |
  Catharine
- |
  catharses
- |
  catharsis
- |
  cathartic
- |
  Cathay
- |
  cathectic
- |
  cathedral
- |
  Cather
- |
  Catherine
- |
  catheter
- |
  catheterize
- |
  cathexis
- |
  Cathie
- |
  Cathleen
- |
  cathodal
- |
  cathode
- |
  cathodic
- |
  Catholic
- |
  catholic
- |
  catholically
- |
  Catholicism
- |
  catholicity
- |
  catholicly
- |
  Cathryn
- |
  Cathy
- |
  Catiline
- |
  cation
- |
  cationic
- |
  catkin
- |
  catlike
- |
  catnap
- |
  catnip
- |
  Catskill
- |
  Catskills
- |
  catspaw
- |
  catsup
- |
  cattail
- |
  cattily
- |
  cattiness
- |
  cattle
- |
  cattleman
- |
  catty
- |
  Catullus
- |
  catwalk
- |
  Caucasia
- |
  Caucasian
- |
  Caucasoid
- |
  Caucasus
- |
  caucus
- |
  caudal
- |
  caudally
- |
  caudillo
- |
  caught
- |
  cauldron
- |
  cauliflower
- |
  caulk
- |
  caulker
- |
  caulking
- |
  causal
- |
  causality
- |
  causally
- |
  causation
- |
  causative
- |
  cause
- |
  causeless
- |
  causer
- |
  causerie
- |
  causeway
- |
  caustic
- |
  caustically
- |
  causticity
- |
  cauterize
- |
  caution
- |
  cautionary
- |
  cautious
- |
  cautiously
- |
  cautiousness
- |
  cavalcade
- |
  Cavalier
- |
  cavalier
- |
  cavalierly
- |
  cavalry
- |
  cavalryman
- |
  caveat
- |
  caveman
- |
  Cavendish
- |
  caver
- |
  cavern
- |
  cavernous
- |
  cavernously
- |
  caviar
- |
  caviare
- |
  cavil
- |
  caviler
- |
  caviller
- |
  caving
- |
  cavitation
- |
  cavity
- |
  cavort
- |
  Cavour
- |
  Caxton
- |
  Cayenne
- |
  cayenne
- |
  Cayman
- |
  cayman
- |
  Cayuga
- |
  Cayuse
- |
  cayuse
- |
  cease
- |
  ceasefire
- |
  ceaseless
- |
  ceaselessly
- |
  Ceausescu
- |
  cecal
- |
  cecally
- |
  Cecelia
- |
  Cecil
- |
  Cecile
- |
  Cecilia
- |
  Cecily
- |
  cecum
- |
  cedar
- |
  ceder
- |
  cedilla
- |
  Cedric
- |
  ceiba
- |
  ceilidh
- |
  ceiling
- |
  celadon
- |
  celandine
- |
  Celebes
- |
  celebrant
- |
  celebrate
- |
  celebrated
- |
  celebration
- |
  celebrator
- |
  celebratory
- |
  celebrity
- |
  celerity
- |
  celery
- |
  celesta
- |
  Celeste
- |
  celeste
- |
  celestial
- |
  celestially
- |
  Celia
- |
  celibacy
- |
  celibate
- |
  cellar
- |
  cellaret
- |
  cellarette
- |
  cellblock
- |
  celled
- |
  celli
- |
  Cellini
- |
  cellist
- |
  cellmate
- |
  cello
- |
  cellophane
- |
  cellular
- |
  cellularity
- |
  cellulite
- |
  celluloid
- |
  cellulose
- |
  cellulosic
- |
  Celsius
- |
  Celtic
- |
  Celticism
- |
  Celticist
- |
  cembali
- |
  cembalist
- |
  cembalo
- |
  cement
- |
  cementer
- |
  cementum
- |
  cemetery
- |
  cenacle
- |
  cenobite
- |
  cenobitic
- |
  cenobitical
- |
  cenotaph
- |
  Cenozoic
- |
  censer
- |
  censor
- |
  censorial
- |
  censorious
- |
  censoriously
- |
  censorship
- |
  censurable
- |
  censure
- |
  censurer
- |
  census
- |
  centaur
- |
  Centaurus
- |
  centavo
- |
  centenarian
- |
  centenary
- |
  centennial
- |
  center
- |
  centerboard
- |
  centered
- |
  centerfold
- |
  centerpiece
- |
  centesimal
- |
  centesimally
- |
  centesimo
- |
  Centigrade
- |
  centigrade
- |
  centigram
- |
  centiliter
- |
  centime
- |
  centimeter
- |
  centimetre
- |
  centimo
- |
  centipede
- |
  Central
- |
  central
- |
  centralise
- |
  centrality
- |
  centralize
- |
  centralizer
- |
  centrally
- |
  centre
- |
  centred
- |
  centrepiece
- |
  centrifugal
- |
  centrifuge
- |
  centripetal
- |
  centrism
- |
  centrist
- |
  centurion
- |
  century
- |
  cephalic
- |
  cephalopod
- |
  Cepheus
- |
  ceramic
- |
  ceramicist
- |
  ceramics
- |
  ceramist
- |
  Cerberus
- |
  cereal
- |
  cerebella
- |
  cerebellar
- |
  cerebellum
- |
  cerebra
- |
  cerebral
- |
  cerebrally
- |
  cerebrate
- |
  cerebration
- |
  cerebrum
- |
  cerecloth
- |
  cerement
- |
  cerements
- |
  ceremonial
- |
  ceremonially
- |
  ceremonious
- |
  ceremony
- |
  Ceres
- |
  cereus
- |
  cerise
- |
  cerium
- |
  cermet
- |
  certain
- |
  certainly
- |
  certainty
- |
  certifiable
- |
  certifiably
- |
  certificate
- |
  certified
- |
  certifier
- |
  certify
- |
  certitude
- |
  cerulean
- |
  cerumen
- |
  ceruminous
- |
  Cervantes
- |
  cervical
- |
  cervices
- |
  cervine
- |
  cervix
- |
  Cesarean
- |
  cesarean
- |
  Cesarian
- |
  cesarian
- |
  cesium
- |
  cessation
- |
  cession
- |
  cesspool
- |
  cesura
- |
  cesurae
- |
  cetacean
- |
  cetaceous
- |
  Cetus
- |
  Ceuta
- |
  Ceylon
- |
  Ceylonese
- |
  Cezanne
- |
  Chablis
- |
  chadar
- |
  Chadian
- |
  Chadic
- |
  chador
- |
  chafe
- |
  chafer
- |
  chaff
- |
  chaffer
- |
  chafferer
- |
  chaffinch
- |
  chaffy
- |
  Chagall
- |
  Chagos
- |
  chagrin
- |
  chain
- |
  chained
- |
  chains
- |
  chainsaw
- |
  chair
- |
  chairlift
- |
  chairman
- |
  chairmanship
- |
  chairperson
- |
  chairwoman
- |
  chaise
- |
  chalcedonic
- |
  chalcedony
- |
  chalcopyrite
- |
  Chaldaea
- |
  Chaldea
- |
  Chaldean
- |
  Chaldee
- |
  chalet
- |
  chalice
- |
  chalk
- |
  chalkboard
- |
  chalkiness
- |
  chalky
- |
  challah
- |
  challenge
- |
  challenged
- |
  challenger
- |
  challenging
- |
  challie
- |
  challis
- |
  challot
- |
  challoth
- |
  Chamaeleon
- |
  chamaeleon
- |
  chamber
- |
  chambered
- |
  Chamberlain
- |
  chamberlain
- |
  chambermaid
- |
  chambers
- |
  chambray
- |
  chameleon
- |
  chameleonic
- |
  chamfer
- |
  chammy
- |
  chamois
- |
  chamoix
- |
  chamomile
- |
  champ
- |
  Champagne
- |
  champagne
- |
  Champaign
- |
  champaign
- |
  champion
- |
  championship
- |
  Champlain
- |
  chance
- |
  chancel
- |
  chancellery
- |
  Chancellor
- |
  chancellor
- |
  chancellory
- |
  chancery
- |
  chances
- |
  chanciness
- |
  chancre
- |
  chancroid
- |
  chancrous
- |
  chancy
- |
  chandelier
- |
  Chandigarh
- |
  Chandler
- |
  chandler
- |
  chandlery
- |
  Chanel
- |
  Chang
- |
  Changchun
- |
  change
- |
  changeable
- |
  changeful
- |
  changeless
- |
  changeling
- |
  changeover
- |
  changer
- |
  Changsha
- |
  channel
- |
  channelize
- |
  channels
- |
  chanson
- |
  chant
- |
  chanter
- |
  chanteuse
- |
  chantey
- |
  chanticleer
- |
  chanting
- |
  chanty
- |
  Chanukah
- |
  Chaos
- |
  chaos
- |
  chaotic
- |
  chaotically
- |
  chaparral
- |
  chapati
- |
  chapbook
- |
  chapeau
- |
  chapeaux
- |
  chapel
- |
  chaperon
- |
  chaperonage
- |
  chaperone
- |
  chapfallen
- |
  chaplain
- |
  chaplaincy
- |
  chaplainship
- |
  chaplet
- |
  chapleted
- |
  Chaplin
- |
  Chapman
- |
  chapman
- |
  chapped
- |
  chaps
- |
  chapter
- |
  character
- |
  characterise
- |
  characterize
- |
  charade
- |
  charades
- |
  charbroil
- |
  charcoal
- |
  chard
- |
  chardonnay
- |
  charge
- |
  chargeable
- |
  charged
- |
  charger
- |
  charily
- |
  chariness
- |
  chariot
- |
  charioteer
- |
  charisma
- |
  charismata
- |
  charismatic
- |
  charitable
- |
  charitably
- |
  Charity
- |
  charity
- |
  charivari
- |
  charlatan
- |
  charlatanism
- |
  charlatanry
- |
  Charlemagne
- |
  Charlene
- |
  Charleroi
- |
  Charles
- |
  Charleston
- |
  Charlotte
- |
  charm
- |
  charmed
- |
  charmer
- |
  charming
- |
  charmingly
- |
  charmless
- |
  charnel
- |
  Charon
- |
  charred
- |
  charring
- |
  chart
- |
  charter
- |
  chartered
- |
  charterer
- |
  Chartres
- |
  chartreuse
- |
  charwoman
- |
  chary
- |
  Charybdis
- |
  Chase
- |
  chase
- |
  chaser
- |
  Chasid
- |
  Chasidim
- |
  chasm
- |
  chasmic
- |
  chasse
- |
  Chassid
- |
  Chassidic
- |
  Chassidim
- |
  Chassidism
- |
  chassis
- |
  chaste
- |
  chastely
- |
  chasten
- |
  chastener
- |
  chasteness
- |
  chastise
- |
  chastisement
- |
  chastiser
- |
  chastity
- |
  chasuble
- |
  chateau
- |
  chateaux
- |
  chatelaine
- |
  chatoyance
- |
  chatoyancy
- |
  chatoyant
- |
  chatroom
- |
  Chattanooga
- |
  chattel
- |
  chatter
- |
  chatterbox
- |
  chatterer
- |
  Chatterton
- |
  chattily
- |
  chattiness
- |
  chatty
- |
  Chaucer
- |
  Chaucerian
- |
  chauffeur
- |
  Chauncey
- |
  chaunt
- |
  Chautauqua
- |
  chautauqua
- |
  chauvinism
- |
  chauvinist
- |
  chauvinistic
- |
  Chavez
- |
  cheap
- |
  cheapen
- |
  cheaply
- |
  cheapness
- |
  cheapskate
- |
  cheat
- |
  cheater
- |
  cheating
- |
  cheatingly
- |
  Cheboksary
- |
  Chechen
- |
  Chechnya
- |
  check
- |
  checkable
- |
  checkbook
- |
  checked
- |
  checker
- |
  checkerberry
- |
  checkerboard
- |
  checkered
- |
  checkers
- |
  checklist
- |
  checkmate
- |
  checkoff
- |
  checkout
- |
  checkpoint
- |
  checkrein
- |
  checkroom
- |
  checkup
- |
  Cheddar
- |
  cheddar
- |
  cheek
- |
  cheekbone
- |
  cheeked
- |
  cheekily
- |
  cheekiness
- |
  cheeky
- |
  cheep
- |
  cheeper
- |
  cheer
- |
  cheerer
- |
  cheerful
- |
  cheerfully
- |
  cheerfulness
- |
  cheerily
- |
  cheeriness
- |
  cheering
- |
  cheerio
- |
  cheerleader
- |
  cheerless
- |
  cheerlessly
- |
  cheers
- |
  cheery
- |
  cheese
- |
  cheeseburger
- |
  cheesecake
- |
  cheesecloth
- |
  cheeseparing
- |
  cheesiness
- |
  cheesy
- |
  cheetah
- |
  Cheever
- |
  Chekhov
- |
  Chekhovian
- |
  Chelmsford
- |
  Chelyabinsk
- |
  chemical
- |
  chemically
- |
  chemise
- |
  chemist
- |
  chemistry
- |
  Chemnitz
- |
  chemo
- |
  chemotherapy
- |
  chemurgic
- |
  chemurgical
- |
  chemurgy
- |
  Chengchou
- |
  Chengchow
- |
  Chengdu
- |
  Chengtu
- |
  chenille
- |
  Chennai
- |
  Cheops
- |
  cheque
- |
  chequer
- |
  Cherepovets
- |
  Cherie
- |
  cherish
- |
  cherishable
- |
  cherished
- |
  cherisher
- |
  Chernenko
- |
  Chernobyl
- |
  chernozem
- |
  Cherokee
- |
  cheroot
- |
  Cherry
- |
  cherry
- |
  cherrystone
- |
  chert
- |
  cherty
- |
  cherub
- |
  cherubic
- |
  cherubically
- |
  cherubim
- |
  chervil
- |
  Cheryl
- |
  Chesapeake
- |
  Cheshire
- |
  chess
- |
  chessboard
- |
  chessman
- |
  chest
- |
  chested
- |
  Chester
- |
  Chesterfield
- |
  chesterfield
- |
  Chesterton
- |
  chestful
- |
  chestily
- |
  chestiness
- |
  chestnut
- |
  chesty
- |
  chetrum
- |
  Chetumal
- |
  Chevalier
- |
  chevalier
- |
  Cheviot
- |
  cheviot
- |
  chevre
- |
  chevron
- |
  chewable
- |
  chewer
- |
  chewiness
- |
  chewy
- |
  Cheyenne
- |
  Chiai
- |
  Chianti
- |
  Chiapas
- |
  chiaroscuro
- |
  chiasmus
- |
  chiastic
- |
  Chiba
- |
  Chicago
- |
  Chicagoan
- |
  Chicana
- |
  chicane
- |
  chicanery
- |
  Chicano
- |
  Chichester
- |
  chichi
- |
  chick
- |
  chickadee
- |
  Chickasaw
- |
  chicken
- |
  chickenfeed
- |
  chickenpox
- |
  chickpea
- |
  chickweed
- |
  Chiclayo
- |
  chicle
- |
  chicly
- |
  chicness
- |
  chicory
- |
  chidden
- |
  chide
- |
  chider
- |
  chidingly
- |
  Chief
- |
  chief
- |
  chiefdom
- |
  chiefly
- |
  chieftain
- |
  chieftaincy
- |
  chiffon
- |
  chiffonier
- |
  Chifley
- |
  chigger
- |
  chignon
- |
  chigoe
- |
  Chihuahua
- |
  chihuahua
- |
  chilblain
- |
  chilblained
- |
  child
- |
  childbearing
- |
  childbirth
- |
  childcare
- |
  childhood
- |
  childish
- |
  childishly
- |
  childishness
- |
  childless
- |
  childlike
- |
  childproof
- |
  children
- |
  Chile
- |
  chile
- |
  Chilean
- |
  chili
- |
  chiliad
- |
  chiliasm
- |
  chiliast
- |
  chiliastic
- |
  chiliburger
- |
  chilidog
- |
  Chilin
- |
  chill
- |
  chiller
- |
  chilli
- |
  chilliness
- |
  chilling
- |
  chillingly
- |
  chillness
- |
  chilly
- |
  Chilpancingo
- |
  Chilung
- |
  chimaera
- |
  Chimborazo
- |
  Chimbote
- |
  chime
- |
  chimer
- |
  Chimera
- |
  chimera
- |
  chimeric
- |
  chimerical
- |
  chimerically
- |
  chimes
- |
  chimney
- |
  chimneypiece
- |
  chimp
- |
  chimpanzee
- |
  China
- |
  china
- |
  Chinan
- |
  Chinatown
- |
  chinaware
- |
  chinch
- |
  chinchilla
- |
  Chinchow
- |
  chine
- |
  Chinese
- |
  chink
- |
  chinless
- |
  chino
- |
  chinoiserie
- |
  Chinook
- |
  chinook
- |
  Chinookan
- |
  chinos
- |
  chinquapin
- |
  chintz
- |
  chintzily
- |
  chintziness
- |
  chintzy
- |
  Chipewayan
- |
  Chipewyan
- |
  chipmunk
- |
  chipped
- |
  chipper
- |
  Chippewa
- |
  chips
- |
  Chirac
- |
  Chirico
- |
  chirographic
- |
  chirography
- |
  chiromancer
- |
  chiromancy
- |
  chiropodist
- |
  chiropody
- |
  chiropractic
- |
  chiropractor
- |
  chirp
- |
  chirrup
- |
  chisel
- |
  chiseled
- |
  chiseler
- |
  chiseller
- |
  Chisinau
- |
  Chita
- |
  chitchat
- |
  chitin
- |
  chitinous
- |
  chitlings
- |
  chitlins
- |
  chiton
- |
  Chittagong
- |
  chitterlings
- |
  chivalric
- |
  chivalrous
- |
  chivalrously
- |
  chivalry
- |
  chive
- |
  chives
- |
  chlamydia
- |
  chlamydiae
- |
  Chloe
- |
  chloral
- |
  chlorate
- |
  chlordan
- |
  chlordane
- |
  chlorella
- |
  chloride
- |
  chloridic
- |
  chlorinate
- |
  chlorination
- |
  chlorinator
- |
  chlorine
- |
  chlorite
- |
  chloroform
- |
  chlorophyll
- |
  chloroplast
- |
  chocaholic
- |
  chock
- |
  chockablock
- |
  chockfull
- |
  chocoholic
- |
  chocolate
- |
  chocolatey
- |
  chocolatier
- |
  chocolaty
- |
  Choctaw
- |
  choice
- |
  choiceness
- |
  choir
- |
  choirboy
- |
  choirmaster
- |
  choke
- |
  choker
- |
  choler
- |
  cholera
- |
  choleraic
- |
  choleric
- |
  cholerically
- |
  cholesterol
- |
  cholla
- |
  chomp
- |
  Chomsky
- |
  Chongjin
- |
  Chongqing
- |
  Chonju
- |
  choose
- |
  chooser
- |
  choosey
- |
  choosiness
- |
  choosy
- |
  chophouse
- |
  Chopin
- |
  chopper
- |
  choppers
- |
  choppily
- |
  choppiness
- |
  choppy
- |
  chops
- |
  chopstick
- |
  chopsticks
- |
  choral
- |
  chorale
- |
  chorally
- |
  chord
- |
  chordal
- |
  chordate
- |
  chore
- |
  chorea
- |
  choregrapher
- |
  choregraphic
- |
  choregraphy
- |
  choreograph
- |
  choreography
- |
  chores
- |
  chorioid
- |
  chorister
- |
  chorizo
- |
  choroid
- |
  chortle
- |
  chortler
- |
  chorus
- |
  chose
- |
  chosen
- |
  chowchow
- |
  chowder
- |
  chrestomathy
- |
  Chretien
- |
  Chris
- |
  chrism
- |
  chrismal
- |
  chrisom
- |
  Christ
- |
  Christchurch
- |
  christen
- |
  Christendom
- |
  christening
- |
  Christian
- |
  christiania
- |
  Christianity
- |
  Christianize
- |
  Christianly
- |
  Christie
- |
  christie
- |
  Christina
- |
  Christine
- |
  Christlike
- |
  Christly
- |
  Christmas
- |
  Christopher
- |
  Christy
- |
  christy
- |
  chromatic
- |
  chromaticism
- |
  chromatin
- |
  chrome
- |
  chromium
- |
  chromosomal
- |
  chromosome
- |
  chromosphere
- |
  chronic
- |
  chronically
- |
  chronicity
- |
  chronicle
- |
  chronicler
- |
  Chronicles
- |
  chronograph
- |
  chronography
- |
  chronologic
- |
  chronologist
- |
  chronology
- |
  chronometer
- |
  chronometric
- |
  chronometry
- |
  chrysalid
- |
  chrysalides
- |
  chrysalis
- |
  chthonian
- |
  chthonic
- |
  chubbily
- |
  chubbiness
- |
  chubby
- |
  chuck
- |
  chuckhole
- |
  chuckle
- |
  chuckwalla
- |
  chuddar
- |
  chugalug
- |
  chukka
- |
  chukkar
- |
  chukker
- |
  Chumash
- |
  chummily
- |
  chumminess
- |
  chummy
- |
  chump
- |
  Chungking
- |
  chunk
- |
  chunkiness
- |
  chunky
- |
  Church
- |
  church
- |
  churchgoer
- |
  churchgoing
- |
  Churchill
- |
  Churchillian
- |
  churchless
- |
  churchman
- |
  churchwarden
- |
  churchwoman
- |
  churchyard
- |
  churl
- |
  churlish
- |
  churlishly
- |
  churlishness
- |
  churn
- |
  churner
- |
  chute
- |
  chutnee
- |
  chutney
- |
  chutzpa
- |
  chutzpah
- |
  chyle
- |
  chylous
- |
  chyme
- |
  chymous
- |
  ciboria
- |
  ciborium
- |
  cicada
- |
  cicadae
- |
  cicatrice
- |
  cicatrices
- |
  cicatricial
- |
  cicatrix
- |
  Cicely
- |
  Cicero
- |
  cicerone
- |
  ciceroni
- |
  Ciceronian
- |
  cider
- |
  cigar
- |
  cigaret
- |
  cigarette
- |
  cigarillo
- |
  cilantro
- |
  cilia
- |
  ciliary
- |
  ciliate
- |
  ciliated
- |
  cilium
- |
  cimetidine
- |
  cinch
- |
  cinchona
- |
  Cincinnati
- |
  Cincinnatus
- |
  cincture
- |
  cinder
- |
  Cinderella
- |
  cinders
- |
  cindery
- |
  Cindy
- |
  cineast
- |
  cineaste
- |
  cinema
- |
  cinematheque
- |
  cinematic
- |
  cinematize
- |
  cineraria
- |
  cinerarium
- |
  cinerary
- |
  cinereous
- |
  cinnabar
- |
  cinnamon
- |
  cinquecento
- |
  cinquefoil
- |
  cioppino
- |
  cipher
- |
  circa
- |
  circadian
- |
  Circe
- |
  Circinus
- |
  circle
- |
  circler
- |
  circlet
- |
  circuit
- |
  circuital
- |
  circuitous
- |
  circuitously
- |
  circuitry
- |
  circuity
- |
  circular
- |
  circularity
- |
  circularize
- |
  circularizer
- |
  circularly
- |
  circulate
- |
  circulation
- |
  circulative
- |
  circulator
- |
  circulatory
- |
  circumcise
- |
  circumcision
- |
  circumflex
- |
  circumlunar
- |
  circumpolar
- |
  circumscribe
- |
  circumsolar
- |
  circumspect
- |
  circumstance
- |
  circumvent
- |
  circus
- |
  circusy
- |
  cirque
- |
  cirrhoses
- |
  cirrhosis
- |
  cirrhotic
- |
  cirri
- |
  cirrocumulus
- |
  cirrostratus
- |
  cirrus
- |
  cislunar
- |
  cistern
- |
  citable
- |
  citadel
- |
  citation
- |
  citification
- |
  citified
- |
  citify
- |
  citizen
- |
  citizenly
- |
  citizenry
- |
  citizenship
- |
  citrate
- |
  citric
- |
  citrine
- |
  citron
- |
  citronella
- |
  citrous
- |
  citrus
- |
  civet
- |
  civic
- |
  civically
- |
  civics
- |
  civies
- |
  civil
- |
  civilian
- |
  civilisation
- |
  civilise
- |
  civilised
- |
  civilities
- |
  civility
- |
  civilization
- |
  civilize
- |
  civilized
- |
  civilizer
- |
  civilly
- |
  civvies
- |
  clabber
- |
  clack
- |
  clacker
- |
  claddagh
- |
  cladding
- |
  cladism
- |
  cladistic
- |
  cladistics
- |
  claim
- |
  claimable
- |
  claimant
- |
  claimer
- |
  clairaudient
- |
  Claire
- |
  clairvoyance
- |
  clairvoyant
- |
  clamant
- |
  clamantly
- |
  clambake
- |
  clamber
- |
  clamberer
- |
  clammer
- |
  clammily
- |
  clamminess
- |
  clammy
- |
  clamor
- |
  clamorous
- |
  clamorously
- |
  clamour
- |
  clamp
- |
  clampdown
- |
  clamper
- |
  clamping
- |
  clamshell
- |
  clandestine
- |
  clang
- |
  clangor
- |
  clangorous
- |
  clangorously
- |
  clangour
- |
  clank
- |
  clannish
- |
  clannishly
- |
  clannishness
- |
  clansman
- |
  clanswoman
- |
  clapboard
- |
  clapper
- |
  clapping
- |
  Clapton
- |
  claptrap
- |
  claque
- |
  Clara
- |
  Clare
- |
  Clarence
- |
  claret
- |
  Clarice
- |
  clarify
- |
  clarinet
- |
  clarinetist
- |
  clarinettist
- |
  clarion
- |
  Clarissa
- |
  clarity
- |
  Clark
- |
  Clarke
- |
  clash
- |
  clasp
- |
  class
- |
  classic
- |
  classical
- |
  classicalism
- |
  classicality
- |
  classically
- |
  classicism
- |
  classicist
- |
  Classics
- |
  classics
- |
  classifiable
- |
  classified
- |
  classifier
- |
  classify
- |
  classily
- |
  classiness
- |
  classism
- |
  classist
- |
  classless
- |
  classmate
- |
  classroom
- |
  classwork
- |
  classy
- |
  clastic
- |
  clatter
- |
  Claud
- |
  Claude
- |
  Claudette
- |
  Claudia
- |
  Claudine
- |
  Claudius
- |
  clausal
- |
  clause
- |
  Clausewitz
- |
  claustral
- |
  clavichord
- |
  clavicle
- |
  clavier
- |
  clawed
- |
  clayey
- |
  clayish
- |
  Claymation
- |
  claymore
- |
  Clayton
- |
  clean
- |
  cleanable
- |
  cleaner
- |
  cleaners
- |
  cleaning
- |
  cleanliness
- |
  cleanly
- |
  cleanness
- |
  cleanse
- |
  cleanser
- |
  cleanup
- |
  clear
- |
  clearance
- |
  clearcut
- |
  clearheaded
- |
  clearing
- |
  clearly
- |
  clearness
- |
  clearstory
- |
  Clearwater
- |
  cleat
- |
  cleats
- |
  cleavable
- |
  cleavage
- |
  cleave
- |
  cleaver
- |
  cleft
- |
  clematis
- |
  Clemenceau
- |
  clemency
- |
  Clemens
- |
  Clement
- |
  clement
- |
  Clementina
- |
  Clementine
- |
  clemently
- |
  clench
- |
  Cleopatra
- |
  clerestory
- |
  clergy
- |
  clergyman
- |
  clergywoman
- |
  cleric
- |
  clerical
- |
  clericalism
- |
  clericalist
- |
  clerically
- |
  clerk
- |
  clerkship
- |
  Cleveland
- |
  clever
- |
  cleverly
- |
  cleverness
- |
  clevis
- |
  cliche
- |
  cliched
- |
  click
- |
  clicker
- |
  client
- |
  clientele
- |
  clientship
- |
  cliff
- |
  cliffhanger
- |
  Clifford
- |
  cliffy
- |
  Clifton
- |
  climacteric
- |
  climactic
- |
  climate
- |
  climatic
- |
  climatical
- |
  climatically
- |
  climatologic
- |
  climatology
- |
  climax
- |
  climb
- |
  climbable
- |
  climber
- |
  climbing
- |
  clime
- |
  climes
- |
  clinch
- |
  clincher
- |
  cling
- |
  clinger
- |
  clinging
- |
  clingstone
- |
  clingy
- |
  clinic
- |
  clinical
- |
  clinically
- |
  clinician
- |
  clink
- |
  clinker
- |
  Clint
- |
  Clinton
- |
  cliometric
- |
  cliometrics
- |
  clipboard
- |
  clipped
- |
  clipper
- |
  clippers
- |
  clipping
- |
  clips
- |
  clique
- |
  cliquey
- |
  cliquish
- |
  cliquishly
- |
  cliquishness
- |
  cliquy
- |
  clitoral
- |
  clitorides
- |
  clitoris
- |
  Clive
- |
  cloaca
- |
  cloacae
- |
  cloak
- |
  cloakroom
- |
  clobber
- |
  cloche
- |
  clock
- |
  clocker
- |
  clockwise
- |
  clockwork
- |
  cloddish
- |
  cloddishly
- |
  cloddishness
- |
  cloddy
- |
  clodhopper
- |
  clodhoppers
- |
  clogged
- |
  cloggy
- |
  clogs
- |
  cloisonne
- |
  cloister
- |
  cloistered
- |
  cloistral
- |
  clomp
- |
  clonal
- |
  clone
- |
  clonk
- |
  closable
- |
  close
- |
  closeable
- |
  closed
- |
  closefisted
- |
  closefitting
- |
  closely
- |
  closemouthed
- |
  closeness
- |
  closeout
- |
  closet
- |
  closeted
- |
  closeup
- |
  closing
- |
  closure
- |
  cloth
- |
  clothe
- |
  clothed
- |
  clothes
- |
  clotheshorse
- |
  clothesline
- |
  clothespin
- |
  clothespress
- |
  clothier
- |
  clothing
- |
  Clotho
- |
  cloture
- |
  cloud
- |
  cloudburst
- |
  cloudily
- |
  cloudiness
- |
  cloudless
- |
  cloudlet
- |
  cloudy
- |
  Clouet
- |
  clout
- |
  clove
- |
  cloven
- |
  clover
- |
  cloverleaf
- |
  cloverleaves
- |
  Clovis
- |
  clown
- |
  clowning
- |
  clownish
- |
  clownishly
- |
  clownishness
- |
  cloying
- |
  cloyingly
- |
  cloyingness
- |
  clubfeet
- |
  clubfoot
- |
  clubfooted
- |
  clubhouse
- |
  cluck
- |
  clueless
- |
  clump
- |
  clumpy
- |
  clumsily
- |
  clumsiness
- |
  clumsy
- |
  clung
- |
  clunk
- |
  clunker
- |
  clunky
- |
  cluster
- |
  clustered
- |
  clutch
- |
  clutches
- |
  clutter
- |
  cluttered
- |
  Clwyd
- |
  Clyde
- |
  Clydesdale
- |
  Clytemnestra
- |
  cnidarian
- |
  coach
- |
  coachman
- |
  coadjutor
- |
  coagulable
- |
  coagulant
- |
  coagulate
- |
  coagulation
- |
  coagulative
- |
  coagulator
- |
  Coahuila
- |
  coalesce
- |
  coalescence
- |
  coalescent
- |
  coalface
- |
  coalition
- |
  coalitional
- |
  coalitionist
- |
  coalmine
- |
  coals
- |
  coarse
- |
  coarsely
- |
  coarsen
- |
  coarseness
- |
  coast
- |
  coastal
- |
  coaster
- |
  coastguard
- |
  coastline
- |
  coated
- |
  coati
- |
  coatimundi
- |
  coating
- |
  coatrack
- |
  coattail
- |
  coauthor
- |
  coaxer
- |
  coaxial
- |
  coaxially
- |
  coaxingly
- |
  cobalt
- |
  cobble
- |
  cobbled
- |
  cobbler
- |
  cobblestone
- |
  Coblenz
- |
  COBOL
- |
  Cobol
- |
  cobra
- |
  cobweb
- |
  cobwebby
- |
  cocain
- |
  cocaine
- |
  cocci
- |
  coccus
- |
  coccygeal
- |
  coccyges
- |
  coccyx
- |
  Cochabamba
- |
  Cochin
- |
  cochineal
- |
  Cochise
- |
  cochlea
- |
  cochleae
- |
  cochlear
- |
  cockade
- |
  cockamamie
- |
  cockamamy
- |
  cockateel
- |
  cockatiel
- |
  cockatoo
- |
  cockatrice
- |
  cockcrow
- |
  cocker
- |
  cockerel
- |
  cockeyed
- |
  cockfight
- |
  cockfighting
- |
  cockily
- |
  cockiness
- |
  cockle
- |
  cockleshell
- |
  Cockney
- |
  cockney
- |
  cockpit
- |
  cockroach
- |
  cockscomb
- |
  cocksure
- |
  cocktail
- |
  cocky
- |
  cocoa
- |
  cocoanut
- |
  coconut
- |
  cocoon
- |
  cocotte
- |
  Cocteau
- |
  coddle
- |
  coddler
- |
  coded
- |
  codein
- |
  codeine
- |
  codependence
- |
  codependency
- |
  codependent
- |
  coder
- |
  codex
- |
  codfish
- |
  codger
- |
  codices
- |
  codicil
- |
  codicillary
- |
  codification
- |
  codifier
- |
  codify
- |
  coding
- |
  codpiece
- |
  coeducation
- |
  coefficient
- |
  coelenterate
- |
  coelom
- |
  coenobite
- |
  coequal
- |
  coequality
- |
  coequally
- |
  coerce
- |
  coercer
- |
  coercible
- |
  coercion
- |
  coercive
- |
  coeternal
- |
  coeternally
- |
  coeternity
- |
  coeval
- |
  coevality
- |
  coevally
- |
  coevolution
- |
  coevolve
- |
  coexist
- |
  coexistence
- |
  coexistent
- |
  coextensive
- |
  coffee
- |
  coffeecake
- |
  coffeehouse
- |
  coffeemaker
- |
  coffeepot
- |
  coffer
- |
  cofferdam
- |
  coffers
- |
  coffin
- |
  cogency
- |
  cogeneration
- |
  cogent
- |
  cogently
- |
  cogitate
- |
  cogitation
- |
  cogitative
- |
  cogitator
- |
  Cognac
- |
  cognac
- |
  cognate
- |
  cognately
- |
  cognateness
- |
  cognition
- |
  cognitional
- |
  cognitive
- |
  cognitively
- |
  cognizable
- |
  cognizance
- |
  cognizant
- |
  cognomen
- |
  cognomina
- |
  cognoscente
- |
  cognoscenti
- |
  cogwheel
- |
  cohabit
- |
  cohabitant
- |
  cohabitation
- |
  cohabiter
- |
  Cohan
- |
  coheir
- |
  cohere
- |
  coherence
- |
  coherency
- |
  coherent
- |
  coherently
- |
  cohesion
- |
  cohesive
- |
  cohesively
- |
  cohesiveness
- |
  cohort
- |
  cohost
- |
  coiffeur
- |
  coiffeuse
- |
  coiffure
- |
  coign
- |
  Coimbatore
- |
  coinage
- |
  coincide
- |
  coincidence
- |
  coincident
- |
  coincidental
- |
  coiner
- |
  coinsurance
- |
  coital
- |
  coition
- |
  coitus
- |
  colander
- |
  Colbert
- |
  coldblooded
- |
  coldly
- |
  coldness
- |
  coldshoulder
- |
  Coleraine
- |
  Coleridge
- |
  Coleridgian
- |
  coleslaw
- |
  Colette
- |
  coleus
- |
  colic
- |
  colicky
- |
  Colima
- |
  Colin
- |
  coliseum
- |
  colitis
- |
  collaborate
- |
  collaborator
- |
  collage
- |
  collagen
- |
  collapse
- |
  collapsible
- |
  collar
- |
  collarbone
- |
  collard
- |
  collards
- |
  collared
- |
  collarless
- |
  collate
- |
  collateral
- |
  collaterally
- |
  collation
- |
  collator
- |
  colleague
- |
  collect
- |
  collectable
- |
  collectanea
- |
  collected
- |
  collectible
- |
  collecting
- |
  collection
- |
  collective
- |
  collectively
- |
  collectivism
- |
  collectivist
- |
  collectivity
- |
  collectivize
- |
  collector
- |
  Colleen
- |
  colleen
- |
  college
- |
  collegia
- |
  collegial
- |
  collegiality
- |
  collegian
- |
  collegiate
- |
  collegium
- |
  collide
- |
  collider
- |
  collie
- |
  collier
- |
  colliery
- |
  collimate
- |
  Collin
- |
  collinear
- |
  collision
- |
  collocate
- |
  collocation
- |
  collodion
- |
  colloid
- |
  colloidal
- |
  colloquia
- |
  colloquial
- |
  colloquially
- |
  colloquium
- |
  colloquy
- |
  collude
- |
  colluder
- |
  collusion
- |
  collusive
- |
  collusively
- |
  Cologne
- |
  cologne
- |
  cologned
- |
  Colombia
- |
  Colombian
- |
  Colombo
- |
  colon
- |
  colone
- |
  Colonel
- |
  colonel
- |
  colonelcy
- |
  colones
- |
  Colonial
- |
  colonial
- |
  colonialism
- |
  colonialist
- |
  colonially
- |
  colonic
- |
  colonise
- |
  colonist
- |
  colonization
- |
  colonize
- |
  colonizer
- |
  colonnade
- |
  colonnaded
- |
  colony
- |
  colophon
- |
  color
- |
  Coloradan
- |
  Colorado
- |
  Coloradoan
- |
  colorant
- |
  coloration
- |
  coloratura
- |
  colorblind
- |
  Colored
- |
  colored
- |
  colorer
- |
  colorfast
- |
  colorfield
- |
  colorful
- |
  colorfully
- |
  colorfulness
- |
  coloring
- |
  colorist
- |
  colorization
- |
  colorize
- |
  colorless
- |
  colorlessly
- |
  colors
- |
  colossal
- |
  colossally
- |
  Colosseum
- |
  colossi
- |
  Colossians
- |
  colossus
- |
  colostomy
- |
  colostrum
- |
  colour
- |
  Coloured
- |
  coloured
- |
  colourful
- |
  colourfully
- |
  colouring
- |
  colourist
- |
  colporteur
- |
  coltish
- |
  coltishly
- |
  coltishness
- |
  Coltrane
- |
  colubrine
- |
  Columba
- |
  columbaria
- |
  columbarium
- |
  Columbia
- |
  columbine
- |
  columbium
- |
  Columbus
- |
  column
- |
  columnar
- |
  columned
- |
  columnist
- |
  comake
- |
  comaker
- |
  Comanche
- |
  comatose
- |
  combat
- |
  combatant
- |
  combative
- |
  combatively
- |
  combed
- |
  comber
- |
  combination
- |
  combine
- |
  combined
- |
  combiner
- |
  combings
- |
  combo
- |
  combust
- |
  combustible
- |
  combustibly
- |
  combustion
- |
  combustive
- |
  comeback
- |
  comedian
- |
  comedic
- |
  comedienne
- |
  comedown
- |
  comedy
- |
  comeliness
- |
  comely
- |
  comer
- |
  comestible
- |
  comestibles
- |
  comet
- |
  comeuppance
- |
  comfit
- |
  comfort
- |
  comfortable
- |
  comfortably
- |
  comforter
- |
  comforting
- |
  comfortingly
- |
  comfrey
- |
  comfy
- |
  comic
- |
  comical
- |
  comicality
- |
  comically
- |
  comicalness
- |
  comics
- |
  coming
- |
  comity
- |
  comma
- |
  command
- |
  commandant
- |
  commandeer
- |
  Commander
- |
  commander
- |
  commanding
- |
  commandment
- |
  commando
- |
  commemorate
- |
  commemorator
- |
  commence
- |
  commencement
- |
  commend
- |
  commendable
- |
  commendably
- |
  commendation
- |
  commendatory
- |
  commender
- |
  commensal
- |
  commensalism
- |
  commensality
- |
  commensurate
- |
  comment
- |
  commentary
- |
  commentate
- |
  commentator
- |
  commerce
- |
  commercial
- |
  commercially
- |
  commie
- |
  commination
- |
  comminatory
- |
  commingle
- |
  commingler
- |
  commiserate
- |
  commiserator
- |
  commissar
- |
  commissarial
- |
  commissariat
- |
  commissary
- |
  commission
- |
  commissioner
- |
  commit
- |
  commitment
- |
  committable
- |
  committal
- |
  committed
- |
  committee
- |
  committeeman
- |
  commode
- |
  commodify
- |
  commodious
- |
  commodiously
- |
  commodity
- |
  Commodore
- |
  commodore
- |
  Commodus
- |
  common
- |
  commonality
- |
  commonalty
- |
  commoner
- |
  commonly
- |
  commonness
- |
  commonplace
- |
  Commons
- |
  commons
- |
  commonsense
- |
  commonweal
- |
  Commonwealth
- |
  commonwealth
- |
  commotion
- |
  communal
- |
  communality
- |
  communalize
- |
  communally
- |
  commune
- |
  communicable
- |
  communicably
- |
  communicant
- |
  communicate
- |
  communicator
- |
  Communion
- |
  communion
- |
  communique
- |
  Communism
- |
  communism
- |
  Communist
- |
  communist
- |
  communistic
- |
  community
- |
  communize
- |
  commutable
- |
  commutation
- |
  commutative
- |
  commutator
- |
  commute
- |
  commuter
- |
  Comoran
- |
  Comorian
- |
  Comoro
- |
  Comoros
- |
  compact
- |
  compacted
- |
  compacter
- |
  compaction
- |
  compactly
- |
  compactness
- |
  compactor
- |
  compadre
- |
  companion
- |
  companionway
- |
  company
- |
  comparable
- |
  comparably
- |
  comparative
- |
  compare
- |
  compared
- |
  comparer
- |
  comparison
- |
  compartment
- |
  compass
- |
  compassion
- |
  compatible
- |
  compatibly
- |
  compatriot
- |
  compeer
- |
  compel
- |
  compelling
- |
  compellingly
- |
  compendia
- |
  compendious
- |
  compendium
- |
  compensate
- |
  compensation
- |
  compensatory
- |
  compete
- |
  competence
- |
  competency
- |
  competent
- |
  competently
- |
  competing
- |
  competition
- |
  competitive
- |
  competitor
- |
  compilation
- |
  compile
- |
  compiler
- |
  complacence
- |
  complacency
- |
  complacent
- |
  complacently
- |
  complain
- |
  complainant
- |
  complainer
- |
  complaint
- |
  complaisance
- |
  complaisant
- |
  compleat
- |
  complected
- |
  complement
- |
  complemental
- |
  complete
- |
  completely
- |
  completeness
- |
  completion
- |
  complex
- |
  complexation
- |
  complexion
- |
  complexional
- |
  complexioned
- |
  complexities
- |
  complexity
- |
  complexly
- |
  complexness
- |
  compliance
- |
  compliancy
- |
  compliant
- |
  compliantly
- |
  complicate
- |
  complicated
- |
  complication
- |
  complicit
- |
  complicity
- |
  compliment
- |
  compliments
- |
  comply
- |
  component
- |
  componential
- |
  comport
- |
  comportment
- |
  compose
- |
  composed
- |
  composedly
- |
  composer
- |
  Composite
- |
  composite
- |
  compositely
- |
  composition
- |
  compositor
- |
  compost
- |
  composting
- |
  composure
- |
  compote
- |
  compound
- |
  compoundable
- |
  compounded
- |
  compounder
- |
  comprehend
- |
  compress
- |
  compressed
- |
  compressible
- |
  compression
- |
  compressive
- |
  compressor
- |
  comprisable
- |
  comprise
- |
  compromise
- |
  compromiser
- |
  compromising
- |
  comptroller
- |
  compulsion
- |
  compulsive
- |
  compulsively
- |
  compulsorily
- |
  compulsory
- |
  compunction
- |
  compunctious
- |
  computable
- |
  computation
- |
  compute
- |
  computer
- |
  computerise
- |
  computerised
- |
  computerize
- |
  computerized
- |
  computing
- |
  comrade
- |
  comradely
- |
  comradeship
- |
  Comsat
- |
  Comte
- |
  Conakry
- |
  conation
- |
  conative
- |
  concatenate
- |
  concave
- |
  concavely
- |
  concaveness
- |
  concavity
- |
  conceal
- |
  concealable
- |
  concealer
- |
  concealment
- |
  concede
- |
  conceder
- |
  conceit
- |
  conceited
- |
  conceitedly
- |
  conceivable
- |
  conceivably
- |
  conceive
- |
  conceiver
- |
  concelebrant
- |
  concelebrate
- |
  concentrate
- |
  concentrated
- |
  concentrator
- |
  concentric
- |
  concentrical
- |
  Concepcion
- |
  concept
- |
  conception
- |
  conceptional
- |
  conceptual
- |
  conceptually
- |
  concern
- |
  concerned
- |
  concerning
- |
  concernment
- |
  concert
- |
  concerted
- |
  concertedly
- |
  concerti
- |
  concertina
- |
  concertinaed
- |
  concertize
- |
  concerto
- |
  concession
- |
  concessional
- |
  concessioner
- |
  conch
- |
  concierge
- |
  conciliar
- |
  conciliate
- |
  conciliation
- |
  conciliative
- |
  conciliator
- |
  conciliatory
- |
  concise
- |
  concisely
- |
  conciseness
- |
  concision
- |
  conclave
- |
  conclude
- |
  concluding
- |
  conclusion
- |
  conclusive
- |
  conclusively
- |
  concoct
- |
  concocter
- |
  concoction
- |
  concoctor
- |
  concomitance
- |
  concomitant
- |
  Concord
- |
  concord
- |
  concordance
- |
  concordanced
- |
  concordant
- |
  concordantly
- |
  concordat
- |
  concourse
- |
  concrescence
- |
  concrescent
- |
  concrete
- |
  concretely
- |
  concreteness
- |
  concretion
- |
  concubinage
- |
  concubinary
- |
  concubine
- |
  concupiscent
- |
  concur
- |
  concurrence
- |
  concurrency
- |
  concurrent
- |
  concurrently
- |
  concurring
- |
  concussion
- |
  concussive
- |
  condemn
- |
  condemnable
- |
  condemnation
- |
  condemnatory
- |
  condemned
- |
  condemner
- |
  condensable
- |
  condensate
- |
  condensation
- |
  condense
- |
  condensed
- |
  condenser
- |
  condensible
- |
  condescend
- |
  condign
- |
  condignly
- |
  condiment
- |
  condition
- |
  conditional
- |
  conditioned
- |
  conditioner
- |
  conditioning
- |
  conditions
- |
  condo
- |
  condole
- |
  condolence
- |
  condom
- |
  condominia
- |
  condominium
- |
  condonable
- |
  condonation
- |
  condone
- |
  condoner
- |
  condor
- |
  Condorcet
- |
  conduce
- |
  conducive
- |
  conduct
- |
  conductance
- |
  conductible
- |
  conduction
- |
  conductive
- |
  conductively
- |
  conductivity
- |
  conductor
- |
  conduit
- |
  condylar
- |
  condyle
- |
  coneflower
- |
  coney
- |
  confab
- |
  confabulate
- |
  confection
- |
  confectioner
- |
  Confederacy
- |
  confederacy
- |
  Confederate
- |
  confederate
- |
  confer
- |
  conferee
- |
  conference
- |
  conferer
- |
  conferment
- |
  conferrable
- |
  conferral
- |
  conferrer
- |
  confess
- |
  confessed
- |
  confessedly
- |
  confession
- |
  confessional
- |
  confessor
- |
  confetti
- |
  confidant
- |
  confidante
- |
  confide
- |
  confidence
- |
  confident
- |
  confidential
- |
  confidently
- |
  confider
- |
  configurable
- |
  configure
- |
  confinable
- |
  confine
- |
  confineable
- |
  confined
- |
  confinement
- |
  confiner
- |
  confines
- |
  confirm
- |
  confirmable
- |
  confirmation
- |
  confirmatory
- |
  confirmed
- |
  confirmedly
- |
  confiscate
- |
  confiscated
- |
  confiscation
- |
  confiscator
- |
  confiscatory
- |
  conflate
- |
  conflation
- |
  conflict
- |
  conflicted
- |
  conflictive
- |
  confluence
- |
  confluent
- |
  conflux
- |
  conform
- |
  conformable
- |
  conformably
- |
  conformance
- |
  conformation
- |
  conformer
- |
  conformism
- |
  conformist
- |
  conformity
- |
  confound
- |
  confounded
- |
  confoundedly
- |
  confounder
- |
  confrere
- |
  confront
- |
  Confucian
- |
  Confucianism
- |
  Confucianist
- |
  Confucius
- |
  confuse
- |
  confused
- |
  confusedly
- |
  confusedness
- |
  confusing
- |
  confusingly
- |
  confusion
- |
  confutable
- |
  confutation
- |
  confute
- |
  confuter
- |
  conga
- |
  congeal
- |
  congealable
- |
  congealed
- |
  congealment
- |
  congelable
- |
  congelation
- |
  congener
- |
  congeneric
- |
  congenial
- |
  congeniality
- |
  congenially
- |
  congenital
- |
  congenitally
- |
  conger
- |
  congeries
- |
  congest
- |
  congested
- |
  congestion
- |
  congestive
- |
  conglomerate
- |
  Congo
- |
  Congolese
- |
  congrats
- |
  congratulate
- |
  congregant
- |
  congregate
- |
  congregation
- |
  congregator
- |
  Congress
- |
  congress
- |
  congressman
- |
  Congreve
- |
  congruence
- |
  congruency
- |
  congruent
- |
  congruently
- |
  congruity
- |
  congruous
- |
  congruously
- |
  conic
- |
  conical
- |
  conically
- |
  conifer
- |
  coniferous
- |
  conjectural
- |
  conjecture
- |
  conjecturer
- |
  conjoin
- |
  conjoiner
- |
  conjoint
- |
  conjointly
- |
  conjugacy
- |
  conjugal
- |
  conjugality
- |
  conjugally
- |
  conjugate
- |
  conjugately
- |
  conjugation
- |
  conjugative
- |
  conjunct
- |
  conjunction
- |
  conjunctiva
- |
  conjunctivae
- |
  conjunctival
- |
  conjunctive
- |
  conjunctly
- |
  conjuncture
- |
  conjuration
- |
  conjure
- |
  conjurer
- |
  conjuror
- |
  conman
- |
  Connacht
- |
  connate
- |
  connatural
- |
  connaturally
- |
  connect
- |
  connectable
- |
  connected
- |
  connecter
- |
  Connecticut
- |
  connection
- |
  connections
- |
  connective
- |
  connectively
- |
  connectivity
- |
  connector
- |
  Connery
- |
  connexion
- |
  Connie
- |
  conniption
- |
  conniptions
- |
  connivance
- |
  connive
- |
  conniver
- |
  connivery
- |
  conniving
- |
  connoisseur
- |
  Connors
- |
  connotation
- |
  connotative
- |
  connote
- |
  connubial
- |
  connubiality
- |
  connubially
- |
  conquer
- |
  conquerable
- |
  conquerer
- |
  conqueror
- |
  conquest
- |
  conquistador
- |
  Conrad
- |
  Conrail
- |
  consanguine
- |
  conscience
- |
  conscious
- |
  consciously
- |
  conscript
- |
  conscription
- |
  consecrate
- |
  consecrated
- |
  consecration
- |
  consecrative
- |
  consecrator
- |
  consecratory
- |
  consecutive
- |
  consensual
- |
  consensually
- |
  consensus
- |
  consent
- |
  consequence
- |
  consequent
- |
  consequently
- |
  conservable
- |
  conservancy
- |
  conservation
- |
  conservatism
- |
  Conservative
- |
  conservative
- |
  conservator
- |
  conservatory
- |
  conserve
- |
  consider
- |
  considerable
- |
  considerably
- |
  considerate
- |
  considered
- |
  considering
- |
  consign
- |
  consignable
- |
  consignee
- |
  consigner
- |
  consignment
- |
  consignor
- |
  consist
- |
  consistence
- |
  consistency
- |
  consistent
- |
  consistently
- |
  consistory
- |
  consolable
- |
  consolation
- |
  consolatory
- |
  console
- |
  consoler
- |
  consolidate
- |
  consolidator
- |
  consoling
- |
  consolingly
- |
  consomme
- |
  consonance
- |
  consonant
- |
  consonantal
- |
  consonantly
- |
  consort
- |
  consortia
- |
  consortium
- |
  conspectus
- |
  conspicuity
- |
  conspicuous
- |
  conspiracy
- |
  conspirator
- |
  conspire
- |
  Constable
- |
  constable
- |
  constabulary
- |
  Constance
- |
  constancy
- |
  constant
- |
  Constanta
- |
  Constantine
- |
  constantly
- |
  constipate
- |
  constipated
- |
  constipation
- |
  constituency
- |
  constituent
- |
  constitute
- |
  Constitution
- |
  constitution
- |
  constitutive
- |
  constrain
- |
  constrained
- |
  constrainer
- |
  constraint
- |
  constrict
- |
  constricted
- |
  constriction
- |
  constrictive
- |
  constrictor
- |
  construable
- |
  construal
- |
  construct
- |
  constructer
- |
  construction
- |
  constructive
- |
  constructor
- |
  construe
- |
  consuetude
- |
  consul
- |
  consular
- |
  consulate
- |
  consulship
- |
  consult
- |
  consultancy
- |
  consultant
- |
  consultation
- |
  consultative
- |
  consumable
- |
  consume
- |
  consumer
- |
  consumerism
- |
  consumerist
- |
  consuming
- |
  consummate
- |
  consummately
- |
  consummation
- |
  consummator
- |
  consumption
- |
  consumptive
- |
  contact
- |
  contagion
- |
  contagious
- |
  contagiously
- |
  contain
- |
  containable
- |
  container
- |
  containerize
- |
  containment
- |
  contaminant
- |
  contaminate
- |
  contaminated
- |
  contaminator
- |
  conte
- |
  contemn
- |
  contemner
- |
  contemnible
- |
  contemnor
- |
  contemplate
- |
  contemplator
- |
  contemporary
- |
  contempt
- |
  contemptible
- |
  contemptibly
- |
  contemptuous
- |
  contend
- |
  contender
- |
  contending
- |
  content
- |
  contented
- |
  contentedly
- |
  contention
- |
  contentious
- |
  contently
- |
  contentment
- |
  contents
- |
  conterminous
- |
  contest
- |
  contestable
- |
  contestant
- |
  contestation
- |
  contester
- |
  context
- |
  contextless
- |
  contextual
- |
  contextually
- |
  contiguity
- |
  contiguous
- |
  contiguously
- |
  continence
- |
  Continent
- |
  continent
- |
  Continental
- |
  continental
- |
  continently
- |
  contingency
- |
  contingent
- |
  contingently
- |
  continua
- |
  continual
- |
  continually
- |
  continuance
- |
  continuation
- |
  continue
- |
  continuer
- |
  continuity
- |
  continuo
- |
  continuous
- |
  continuously
- |
  continuum
- |
  contort
- |
  contorted
- |
  contortion
- |
  contortive
- |
  contour
- |
  contours
- |
  contra
- |
  contraband
- |
  contrabass
- |
  contract
- |
  contractable
- |
  contractible
- |
  contractile
- |
  contraction
- |
  contractions
- |
  contractor
- |
  contractual
- |
  contradance
- |
  contradict
- |
  contradicter
- |
  contradictor
- |
  contrail
- |
  contralto
- |
  contraption
- |
  contrapuntal
- |
  contrarian
- |
  contrariety
- |
  contrarily
- |
  contrariness
- |
  contrariwise
- |
  contrary
- |
  contrast
- |
  contrastable
- |
  contrasting
- |
  contravene
- |
  contravener
- |
  contredanse
- |
  contretemps
- |
  contribute
- |
  contribution
- |
  contributive
- |
  contributor
- |
  contributory
- |
  contrite
- |
  contritely
- |
  contriteness
- |
  contrition
- |
  contrivance
- |
  contrive
- |
  contrived
- |
  contrivedly
- |
  contriver
- |
  control
- |
  controllable
- |
  controllably
- |
  controlled
- |
  controller
- |
  controls
- |
  controversy
- |
  controvert
- |
  contumacious
- |
  contumacy
- |
  contumelious
- |
  contumely
- |
  contuse
- |
  contusion
- |
  conundrum
- |
  conurbation
- |
  convalesce
- |
  convalescent
- |
  convect
- |
  convection
- |
  convectional
- |
  convective
- |
  convenable
- |
  convenance
- |
  convenances
- |
  convene
- |
  convener
- |
  convenience
- |
  convenient
- |
  conveniently
- |
  convenor
- |
  convent
- |
  conventicle
- |
  convention
- |
  conventional
- |
  conventual
- |
  converge
- |
  convergence
- |
  convergency
- |
  convergent
- |
  conversance
- |
  conversancy
- |
  conversant
- |
  conversantly
- |
  conversation
- |
  converse
- |
  conversely
- |
  conversion
- |
  convert
- |
  converter
- |
  convertible
- |
  convertibles
- |
  convertor
- |
  convex
- |
  convexity
- |
  convexly
- |
  convey
- |
  conveyable
- |
  conveyance
- |
  conveyer
- |
  conveyor
- |
  convict
- |
  conviction
- |
  convince
- |
  convinced
- |
  convincing
- |
  convincingly
- |
  convivial
- |
  conviviality
- |
  convivially
- |
  convocation
- |
  convoke
- |
  convoluted
- |
  convolutedly
- |
  convolution
- |
  convoy
- |
  convulse
- |
  convulsion
- |
  convulsions
- |
  convulsive
- |
  convulsively
- |
  cookbook
- |
  cooked
- |
  cooker
- |
  cookery
- |
  cookie
- |
  cooking
- |
  cookout
- |
  Cookstown
- |
  cooktop
- |
  cookware
- |
  cooky
- |
  coolant
- |
  cooler
- |
  Coolidge
- |
  coolie
- |
  cooling
- |
  coolly
- |
  coolness
- |
  coonhound
- |
  coonskin
- |
  Cooper
- |
  cooper
- |
  cooperage
- |
  cooperate
- |
  cooperation
- |
  cooperative
- |
  cooperator
- |
  cooption
- |
  cooptive
- |
  coordinate
- |
  coordinated
- |
  coordinately
- |
  coordination
- |
  coordinative
- |
  coordinator
- |
  cootie
- |
  cooties
- |
  copacetic
- |
  copartner
- |
  copasetic
- |
  copay
- |
  copayment
- |
  Copenhagen
- |
  Copernican
- |
  Copernicus
- |
  copier
- |
  copilot
- |
  coping
- |
  copious
- |
  copiously
- |
  copiousness
- |
  Copland
- |
  Copley
- |
  copper
- |
  copperhead
- |
  coppery
- |
  coppice
- |
  coppiced
- |
  Coppola
- |
  copra
- |
  coprocessor
- |
  copse
- |
  copter
- |
  Coptic
- |
  copula
- |
  copular
- |
  copulate
- |
  copulation
- |
  copulative
- |
  copulatively
- |
  copulatory
- |
  copybook
- |
  copyboy
- |
  copycat
- |
  copydesk
- |
  copyedit
- |
  copyeditor
- |
  copying
- |
  copyist
- |
  copyreader
- |
  copyright
- |
  copyrighted
- |
  copywriter
- |
  copywriting
- |
  coquet
- |
  coquetry
- |
  coquette
- |
  coquettish
- |
  coquettishly
- |
  coracle
- |
  Coral
- |
  coral
- |
  corbeil
- |
  corbel
- |
  Corbusier
- |
  cordage
- |
  Corday
- |
  Cordelia
- |
  corder
- |
  cordial
- |
  cordiality
- |
  cordially
- |
  cordillera
- |
  cordilleran
- |
  Cordilleras
- |
  cordite
- |
  cordless
- |
  Cordoba
- |
  cordoba
- |
  cordon
- |
  Cordova
- |
  Cordovan
- |
  cordovan
- |
  cords
- |
  corduroy
- |
  corduroys
- |
  cordwainer
- |
  corer
- |
  corespondent
- |
  Corey
- |
  Corfu
- |
  corgi
- |
  coria
- |
  coriander
- |
  Corinne
- |
  Corinth
- |
  Corinthian
- |
  Corinthians
- |
  Coriolanus
- |
  corium
- |
  corkage
- |
  corked
- |
  corker
- |
  corklike
- |
  corkscrew
- |
  corky
- |
  cormorant
- |
  cornball
- |
  cornbread
- |
  corncob
- |
  corncrib
- |
  cornea
- |
  corneal
- |
  corned
- |
  Corneille
- |
  Cornelia
- |
  Cornelius
- |
  corner
- |
  cornerback
- |
  cornered
- |
  cornerstone
- |
  cornet
- |
  cornetist
- |
  cornflakes
- |
  cornflower
- |
  cornice
- |
  corniced
- |
  corniche
- |
  cornicing
- |
  cornily
- |
  corniness
- |
  Cornish
- |
  Cornishman
- |
  Cornishwoman
- |
  cornmeal
- |
  cornpone
- |
  cornrow
- |
  cornstalk
- |
  cornstarch
- |
  cornucopia
- |
  cornucopian
- |
  Cornwall
- |
  Cornwallis
- |
  corny
- |
  corolla
- |
  corollary
- |
  corona
- |
  Coronado
- |
  coronae
- |
  coronal
- |
  coronary
- |
  coronation
- |
  coroner
- |
  coronet
- |
  coroneted
- |
  Corot
- |
  corpora
- |
  Corporal
- |
  corporal
- |
  corporality
- |
  corporally
- |
  corporate
- |
  corporately
- |
  corporation
- |
  corporatism
- |
  corporatist
- |
  corporative
- |
  corporeal
- |
  corporeality
- |
  corporeally
- |
  corps
- |
  corpse
- |
  corpsman
- |
  corpulence
- |
  corpulency
- |
  corpulent
- |
  corpus
- |
  corpuscle
- |
  corpuscular
- |
  corral
- |
  correct
- |
  correctable
- |
  correctible
- |
  correction
- |
  correctional
- |
  corrections
- |
  correctitude
- |
  corrective
- |
  correctly
- |
  correctness
- |
  Correggio
- |
  Corregidor
- |
  correlate
- |
  correlation
- |
  correlative
- |
  correspond
- |
  corridor
- |
  corrigenda
- |
  corrigendum
- |
  corrigible
- |
  Corrine
- |
  corroborate
- |
  corroborator
- |
  corrode
- |
  corrodible
- |
  corrosible
- |
  corrosion
- |
  corrosive
- |
  corrosively
- |
  corrugate
- |
  corrugated
- |
  corrugation
- |
  corrupt
- |
  corrupter
- |
  corruptible
- |
  corruption
- |
  corruptive
- |
  corruptly
- |
  corruptness
- |
  corruptor
- |
  corsage
- |
  corsair
- |
  corset
- |
  corsetry
- |
  Corsica
- |
  Corsican
- |
  cortege
- |
  Cortes
- |
  cortex
- |
  Cortez
- |
  cortical
- |
  cortices
- |
  cortisone
- |
  corundum
- |
  coruscate
- |
  coruscation
- |
  corvee
- |
  corvette
- |
  Corvus
- |
  corymb
- |
  coryza
- |
  Cosby
- |
  cosecant
- |
  cosign
- |
  cosignatory
- |
  cosigner
- |
  cosily
- |
  cosine
- |
  cosiness
- |
  cosmetic
- |
  cosmetically
- |
  cosmetician
- |
  cosmetics
- |
  cosmetology
- |
  cosmic
- |
  cosmical
- |
  cosmically
- |
  cosmogonic
- |
  cosmogonical
- |
  cosmogonist
- |
  cosmogony
- |
  cosmographer
- |
  cosmography
- |
  cosmologic
- |
  cosmological
- |
  cosmologist
- |
  cosmology
- |
  cosmonaut
- |
  cosmopolis
- |
  cosmopolitan
- |
  cosmopolite
- |
  cosmos
- |
  cosponsor
- |
  Cossack
- |
  cossack
- |
  cosset
- |
  costal
- |
  costar
- |
  costing
- |
  costive
- |
  costliness
- |
  costly
- |
  costs
- |
  costume
- |
  costumer
- |
  cotangent
- |
  coterie
- |
  coterminous
- |
  cotillion
- |
  cotillon
- |
  Cotonou
- |
  Cotswold
- |
  cottage
- |
  cottager
- |
  cottar
- |
  cotter
- |
  cotton
- |
  cottonmouth
- |
  cottonseed
- |
  cottontail
- |
  cottonwood
- |
  cottony
- |
  cotyledon
- |
  cotyledonous
- |
  couch
- |
  couchant
- |
  Coueism
- |
  cougar
- |
  cough
- |
  coughing
- |
  could
- |
  coulee
- |
  couloir
- |
  coulomb
- |
  council
- |
  councillor
- |
  councilman
- |
  councilor
- |
  councilwoman
- |
  counsel
- |
  counseling
- |
  counselling
- |
  counsellor
- |
  Counselor
- |
  counselor
- |
  Count
- |
  count
- |
  countable
- |
  countdown
- |
  countenance
- |
  countenancer
- |
  counter
- |
  counteract
- |
  counterblast
- |
  counterclaim
- |
  counterfeit
- |
  counterman
- |
  countermand
- |
  counterpane
- |
  counterpart
- |
  counterplot
- |
  counterpoint
- |
  counterpoise
- |
  countersank
- |
  countersign
- |
  countersink
- |
  counterspy
- |
  countersunk
- |
  countertenor
- |
  countervail
- |
  countess
- |
  counting
- |
  countless
- |
  countrified
- |
  country
- |
  countryfied
- |
  countryman
- |
  countryside
- |
  countrywoman
- |
  county
- |
  coupe
- |
  Couperin
- |
  couple
- |
  coupler
- |
  couplet
- |
  coupling
- |
  coupon
- |
  courage
- |
  courageous
- |
  courageously
- |
  Courbet
- |
  courgette
- |
  courier
- |
  course
- |
  courser
- |
  court
- |
  courteous
- |
  courteously
- |
  courter
- |
  courtesan
- |
  courtesy
- |
  courtezan
- |
  courthouse
- |
  courtier
- |
  courtliness
- |
  courtly
- |
  Courtney
- |
  courtroom
- |
  courtship
- |
  courtyard
- |
  couscous
- |
  cousin
- |
  Cousteau
- |
  couth
- |
  couture
- |
  couturier
- |
  couvade
- |
  coven
- |
  covenant
- |
  covenantal
- |
  covenanter
- |
  covenantor
- |
  Coventry
- |
  cover
- |
  coverage
- |
  coverall
- |
  coveralls
- |
  covered
- |
  covering
- |
  coverlet
- |
  covers
- |
  covert
- |
  covertly
- |
  covertness
- |
  coverture
- |
  coverup
- |
  covet
- |
  coveted
- |
  covetous
- |
  covetously
- |
  covetousness
- |
  covey
- |
  Coward
- |
  coward
- |
  cowardice
- |
  cowardliness
- |
  cowardly
- |
  cowbird
- |
  cowboy
- |
  cowcatcher
- |
  cower
- |
  cowgirl
- |
  cowhand
- |
  cowherd
- |
  cowhide
- |
  Cowley
- |
  cowlick
- |
  cowling
- |
  cowman
- |
  coworker
- |
  Cowpens
- |
  Cowper
- |
  cowpoke
- |
  cowpox
- |
  cowpuncher
- |
  cowrie
- |
  cowry
- |
  cowslip
- |
  coxcomb
- |
  coxcombry
- |
  coxswain
- |
  coyly
- |
  coyness
- |
  coyote
- |
  coypu
- |
  cozen
- |
  cozenage
- |
  cozener
- |
  cozily
- |
  coziness
- |
  Cozumel
- |
  crabbed
- |
  crabbedly
- |
  crabbedness
- |
  crabbily
- |
  crabbiness
- |
  crabby
- |
  crabgrass
- |
  crablike
- |
  crack
- |
  crackdown
- |
  cracked
- |
  cracker
- |
  crackerjack
- |
  crackers
- |
  cracking
- |
  crackle
- |
  crackly
- |
  crackpot
- |
  crackup
- |
  Cracow
- |
  cradle
- |
  cradleboard
- |
  cradlesong
- |
  craft
- |
  craftily
- |
  craftiness
- |
  craftsman
- |
  craftsperson
- |
  craftswoman
- |
  crafty
- |
  cragginess
- |
  craggy
- |
  Craig
- |
  Craigavon
- |
  Craiova
- |
  crammed
- |
  cramp
- |
  cramped
- |
  cramping
- |
  crampon
- |
  cramps
- |
  Cranach
- |
  cranberry
- |
  Crane
- |
  crane
- |
  crania
- |
  cranial
- |
  craniology
- |
  cranium
- |
  crank
- |
  crankcase
- |
  crankily
- |
  crankiness
- |
  crankshaft
- |
  cranky
- |
  Cranmer
- |
  crannied
- |
  cranny
- |
  crape
- |
  crappie
- |
  crappy
- |
  craps
- |
  crapshoot
- |
  crapshooter
- |
  crapulence
- |
  crapulent
- |
  crapulous
- |
  crapy
- |
  craquelure
- |
  crash
- |
  crass
- |
  crassitude
- |
  crassly
- |
  crassness
- |
  Crassus
- |
  crate
- |
  Crater
- |
  crater
- |
  craton
- |
  cravat
- |
  crave
- |
  craven
- |
  cravenly
- |
  cravenness
- |
  craving
- |
  crawdad
- |
  crawfish
- |
  Crawford
- |
  crawl
- |
  crawler
- |
  crawlspace
- |
  crawly
- |
  crayfish
- |
  crayon
- |
  craze
- |
  crazed
- |
  crazily
- |
  craziness
- |
  crazy
- |
  creak
- |
  creakily
- |
  creakiness
- |
  creaky
- |
  cream
- |
  creamer
- |
  creamery
- |
  creamily
- |
  creaminess
- |
  creamy
- |
  crease
- |
  creased
- |
  creaseless
- |
  creaseproof
- |
  create
- |
  Creation
- |
  creation
- |
  creationism
- |
  creationist
- |
  creative
- |
  creatively
- |
  creativeness
- |
  creativity
- |
  Creator
- |
  creator
- |
  creature
- |
  creaturely
- |
  creche
- |
  credence
- |
  credential
- |
  credentials
- |
  credenza
- |
  credibility
- |
  credible
- |
  credibly
- |
  credit
- |
  creditable
- |
  creditably
- |
  creditor
- |
  credits
- |
  Credo
- |
  credo
- |
  credulity
- |
  credulous
- |
  credulously
- |
  creed
- |
  Creek
- |
  creek
- |
  creel
- |
  creep
- |
  creeper
- |
  creepily
- |
  creepiness
- |
  creeping
- |
  creeps
- |
  creepy
- |
  cremains
- |
  cremate
- |
  cremation
- |
  crematoria
- |
  crematorium
- |
  crematory
- |
  creme
- |
  crenelate
- |
  crenelated
- |
  crenelation
- |
  crenellate
- |
  crenellated
- |
  crenellation
- |
  crenshaw
- |
  crenulate
- |
  crenulated
- |
  Creole
- |
  creole
- |
  creosote
- |
  crepe
- |
  crepey
- |
  crepitant
- |
  crepitate
- |
  crepitation
- |
  crept
- |
  crepuscular
- |
  crescendi
- |
  crescendo
- |
  crescent
- |
  crescentic
- |
  cress
- |
  crest
- |
  crested
- |
  crestfallen
- |
  crestless
- |
  Cretaceous
- |
  cretaceous
- |
  Cretan
- |
  Crete
- |
  cretin
- |
  cretinism
- |
  cretinoid
- |
  cretinous
- |
  cretonne
- |
  crevasse
- |
  crevice
- |
  crewcut
- |
  crewed
- |
  crewel
- |
  crewelwork
- |
  crewman
- |
  crewmate
- |
  cribbage
- |
  cribber
- |
  Crick
- |
  crick
- |
  cricket
- |
  cricketeer
- |
  cricketer
- |
  cricketing
- |
  cried
- |
  crier
- |
  crime
- |
  Crimea
- |
  Crimean
- |
  criminal
- |
  criminalist
- |
  criminality
- |
  criminalize
- |
  criminally
- |
  criminology
- |
  crimp
- |
  crimper
- |
  crimson
- |
  cringe
- |
  cringing
- |
  crinkle
- |
  crinkled
- |
  crinkly
- |
  crinoline
- |
  cripple
- |
  crippled
- |
  crippling
- |
  cripplingly
- |
  crises
- |
  crisis
- |
  crisp
- |
  Crispin
- |
  crispiness
- |
  crisply
- |
  crispness
- |
  crispy
- |
  crisscross
- |
  criteria
- |
  criterial
- |
  criterion
- |
  critic
- |
  critical
- |
  criticality
- |
  critically
- |
  criticalness
- |
  criticise
- |
  criticism
- |
  criticizable
- |
  criticize
- |
  criticizer
- |
  critique
- |
  critter
- |
  croak
- |
  croakily
- |
  croakiness
- |
  croaky
- |
  Croat
- |
  Croatia
- |
  Croatian
- |
  Croce
- |
  crochet
- |
  crocheter
- |
  croci
- |
  crock
- |
  crocked
- |
  crockery
- |
  Crockett
- |
  crocodile
- |
  crocodilian
- |
  crocus
- |
  Croesus
- |
  croissant
- |
  Cromwell
- |
  Cromwellian
- |
  crone
- |
  Cronin
- |
  Cronus
- |
  crony
- |
  cronyism
- |
  crook
- |
  crooked
- |
  crookedly
- |
  crookedness
- |
  crookneck
- |
  croon
- |
  crooner
- |
  cropland
- |
  cropped
- |
  cropper
- |
  croquet
- |
  croquette
- |
  Crosby
- |
  crosier
- |
  cross
- |
  crossbar
- |
  crossbeam
- |
  crossbones
- |
  crossbow
- |
  crossbowman
- |
  crossbred
- |
  crossbreed
- |
  crosscheck
- |
  crosscurrent
- |
  crosscut
- |
  crossfire
- |
  crosshair
- |
  crosshatch
- |
  crossing
- |
  crossly
- |
  crossness
- |
  crossover
- |
  crosspatch
- |
  crosspiece
- |
  crossroad
- |
  crossroads
- |
  crosstown
- |
  crosswalk
- |
  crossways
- |
  crosswind
- |
  crosswise
- |
  crossword
- |
  crotch
- |
  crotchet
- |
  crotchety
- |
  crouch
- |
  croup
- |
  croupier
- |
  croupous
- |
  croupy
- |
  crouton
- |
  crowbar
- |
  crowd
- |
  crowded
- |
  crowdedness
- |
  crowfeet
- |
  crowfoot
- |
  Crown
- |
  crown
- |
  crowned
- |
  crowning
- |
  Croydon
- |
  crozier
- |
  cruces
- |
  crucial
- |
  cruciality
- |
  crucially
- |
  crucible
- |
  crucifix
- |
  Crucifixion
- |
  crucifixion
- |
  cruciform
- |
  crucify
- |
  cruddy
- |
  crude
- |
  crudely
- |
  crudeness
- |
  crudites
- |
  crudity
- |
  cruel
- |
  cruelly
- |
  cruelness
- |
  cruelty
- |
  cruet
- |
  Cruikshank
- |
  cruise
- |
  cruiser
- |
  cruising
- |
  cruller
- |
  crumb
- |
  crumble
- |
  crumbliness
- |
  crumbly
- |
  crumby
- |
  crumminess
- |
  crummy
- |
  crumpet
- |
  crumple
- |
  crumpled
- |
  crumply
- |
  crunch
- |
  crunchiness
- |
  crunchy
- |
  crupper
- |
  Crusade
- |
  crusade
- |
  crusader
- |
  Crusades
- |
  cruse
- |
  crush
- |
  crusher
- |
  crushing
- |
  crust
- |
  crustacean
- |
  crustaceous
- |
  crustal
- |
  crustily
- |
  crustiness
- |
  crusty
- |
  crutch
- |
  cruzado
- |
  cruzeiro
- |
  crybaby
- |
  cryer
- |
  crying
- |
  cryogen
- |
  cryogenic
- |
  cryogenics
- |
  cryolite
- |
  cryonic
- |
  cryonics
- |
  cryosurgery
- |
  crypt
- |
  cryptanalyst
- |
  cryptic
- |
  cryptically
- |
  cryptogram
- |
  cryptography
- |
  Crystal
- |
  crystal
- |
  crystalline
- |
  crystallise
- |
  crystallize
- |
  ctenophore
- |
  Cuban
- |
  cubbyhole
- |
  cuber
- |
  cubic
- |
  cubical
- |
  cubically
- |
  cubicle
- |
  cubism
- |
  cubist
- |
  cubistic
- |
  cubit
- |
  cuckold
- |
  cuckoldry
- |
  cuckoo
- |
  cucumber
- |
  Cucuta
- |
  cuddle
- |
  cuddlesome
- |
  cuddly
- |
  cudgel
- |
  Cuenca
- |
  Cuernavaca
- |
  cuesta
- |
  cufflink
- |
  cuffs
- |
  cuirass
- |
  Cuisinart
- |
  cuisine
- |
  Culiacan
- |
  culinarily
- |
  culinary
- |
  Cullen
- |
  culler
- |
  culling
- |
  culminate
- |
  culmination
- |
  culotte
- |
  culottes
- |
  culpability
- |
  culpable
- |
  culpably
- |
  culprit
- |
  cultic
- |
  cultish
- |
  cultism
- |
  cultist
- |
  cultivable
- |
  cultivar
- |
  cultivatable
- |
  cultivate
- |
  cultivated
- |
  cultivation
- |
  cultivator
- |
  cultural
- |
  culturally
- |
  culture
- |
  cultured
- |
  culvert
- |
  cumber
- |
  Cumberland
- |
  cumbersome
- |
  cumbersomely
- |
  Cumbria
- |
  Cumbrian
- |
  cumbrous
- |
  cumbrousness
- |
  cumin
- |
  cummerbund
- |
  Cummings
- |
  cumquat
- |
  cumulative
- |
  cumulatively
- |
  cumuli
- |
  cumulonimbi
- |
  cumulonimbus
- |
  cumulus
- |
  cuneiform
- |
  cunnilinctus
- |
  cunnilingus
- |
  cunning
- |
  cunningly
- |
  Cupar
- |
  cupboard
- |
  cupcake
- |
  cupful
- |
  Cupid
- |
  cupid
- |
  cupidity
- |
  cupola
- |
  cupolaed
- |
  cupreous
- |
  cupric
- |
  curability
- |
  curable
- |
  Curacao
- |
  curacy
- |
  curare
- |
  curari
- |
  curate
- |
  curation
- |
  curative
- |
  curatively
- |
  curator
- |
  curatorial
- |
  curatorship
- |
  curbing
- |
  curbstone
- |
  curdle
- |
  curds
- |
  curdy
- |
  cureless
- |
  curer
- |
  curettage
- |
  curette
- |
  curfew
- |
  Curia
- |
  curia
- |
  Curiae
- |
  curiae
- |
  Curial
- |
  curial
- |
  Curie
- |
  curie
- |
  curio
- |
  curiosa
- |
  curiosity
- |
  curious
- |
  curiously
- |
  curiousness
- |
  Curitiba
- |
  curium
- |
  curler
- |
  curlew
- |
  curlicue
- |
  curliness
- |
  curling
- |
  curly
- |
  curmudgeon
- |
  curmudgeonly
- |
  currant
- |
  currency
- |
  current
- |
  currently
- |
  currentness
- |
  curricula
- |
  curricular
- |
  curriculum
- |
  Currier
- |
  curry
- |
  currycomb
- |
  curse
- |
  cursed
- |
  cursive
- |
  cursively
- |
  cursor
- |
  cursorily
- |
  cursoriness
- |
  cursory
- |
  curst
- |
  curtail
- |
  curtailment
- |
  curtain
- |
  curtal
- |
  Curtin
- |
  Curtis
- |
  Curtiss
- |
  curtly
- |
  curtness
- |
  curtsey
- |
  curtsy
- |
  curvaceous
- |
  curvacious
- |
  curvature
- |
  curve
- |
  curved
- |
  curvet
- |
  curvilinear
- |
  curviness
- |
  curvy
- |
  cushiness
- |
  cushion
- |
  Cushite
- |
  Cushitic
- |
  cushy
- |
  cuspate
- |
  cusped
- |
  cuspid
- |
  cuspidate
- |
  cuspidor
- |
  custard
- |
  Custer
- |
  custodial
- |
  custodian
- |
  custody
- |
  custom
- |
  customarily
- |
  customary
- |
  customer
- |
  customhouse
- |
  customise
- |
  customize
- |
  customs
- |
  cutaneous
- |
  cutaway
- |
  cutback
- |
  cutely
- |
  cuteness
- |
  cutesie
- |
  cutesy
- |
  Cuthbert
- |
  cuticle
- |
  cuticular
- |
  cutlas
- |
  cutlass
- |
  cutler
- |
  cutlery
- |
  cutlet
- |
  cutoff
- |
  cutoffs
- |
  cutout
- |
  cutter
- |
  cutthroat
- |
  cutting
- |
  cuttingly
- |
  cuttlebone
- |
  cuttlefish
- |
  cutup
- |
  cutworm
- |
  Cuvier
- |
  Cuzco
- |
  cyanide
- |
  cyanogen
- |
  cyanosis
- |
  cyanotic
- |
  cybernaut
- |
  cybernetic
- |
  cybernetics
- |
  cyberpunk
- |
  cyberspace
- |
  cyborg
- |
  Cyclades
- |
  cyclamate
- |
  cyclamen
- |
  cycle
- |
  cycler
- |
  cyclic
- |
  cyclical
- |
  cyclically
- |
  cyclicals
- |
  cyclicly
- |
  cycling
- |
  cyclist
- |
  cyclometer
- |
  cyclone
- |
  cyclonic
- |
  cyclopaedia
- |
  cyclopedia
- |
  Cyclopes
- |
  Cyclops
- |
  cyclosporine
- |
  cyclotron
- |
  cyder
- |
  cygnet
- |
  Cygnus
- |
  cylinder
- |
  cylindrical
- |
  cymbal
- |
  cymbalist
- |
  Cymbeline
- |
  Cymric
- |
  Cymru
- |
  Cynic
- |
  cynic
- |
  cynical
- |
  cynically
- |
  cynicism
- |
  cynosure
- |
  Cynthia
- |
  cypher
- |
  cypress
- |
  Cyprian
- |
  Cypriot
- |
  Cypriote
- |
  Cyprus
- |
  Cyrenaic
- |
  Cyrenaica
- |
  Cyrenaican
- |
  Cyrenaicism
- |
  Cyril
- |
  Cyrillic
- |
  Cyrus
- |
  cystic
- |
  cystoscope
- |
  cytologic
- |
  cytological
- |
  cytologist
- |
  cytology
- |
  cytoplasm
- |
  cytoplasmic
- |
  cytosine
- |
  czardom
- |
  czarina
- |
  czarism
- |
  czarist
- |
  Czech
- |
  Czechoslovak
- |
  Czestochowa
- |
  dabber
- |
  dabble
- |
  dabbler
- |
  Dacca
- |
  dacha
- |
  Dachau
- |
  dachshund
- |
  Dacia
- |
  Dacian
- |
  Dacron
- |
  dactyl
- |
  dactylic
- |
  Dadaism
- |
  dadaism
- |
  Dadaist
- |
  dadaist
- |
  Dadaistic
- |
  daddy
- |
  Daedalus
- |
  daemon
- |
  daemonic
- |
  daffily
- |
  daffiness
- |
  daffodil
- |
  daffy
- |
  daftly
- |
  daftness
- |
  dagger
- |
  Dagmar
- |
  daguerrotype
- |
  dahlia
- |
  Dahoman
- |
  Dahomean
- |
  Dahomey
- |
  daikon
- |
  dailiness
- |
  daily
- |
  daimio
- |
  daimon
- |
  daimyo
- |
  daintily
- |
  daintiness
- |
  dainty
- |
  daiquiri
- |
  Dairen
- |
  dairy
- |
  dairying
- |
  dairymaid
- |
  dairyman
- |
  dairywoman
- |
  daishiki
- |
  Daisy
- |
  daisy
- |
  Dakar
- |
  Dakota
- |
  Dakotan
- |
  Dakotas
- |
  dalasi
- |
  Daley
- |
  Dalian
- |
  Daliesque
- |
  Dallas
- |
  Dallasite
- |
  dalliance
- |
  dallier
- |
  dally
- |
  Dalmatia
- |
  Dalmatian
- |
  dalmatian
- |
  Dalton
- |
  damage
- |
  damageable
- |
  damages
- |
  damaging
- |
  Damascene
- |
  damascene
- |
  damascened
- |
  Damascus
- |
  damask
- |
  dammit
- |
  damnable
- |
  damnably
- |
  damnation
- |
  damnatory
- |
  damndest
- |
  damned
- |
  damnedest
- |
  damning
- |
  Damocles
- |
  dampen
- |
  dampener
- |
  damper
- |
  dampish
- |
  damply
- |
  dampness
- |
  damsel
- |
  damselfly
- |
  damson
- |
  Danang
- |
  dance
- |
  danceable
- |
  dancer
- |
  dancing
- |
  dandelion
- |
  dander
- |
  dandify
- |
  dandle
- |
  dandruff
- |
  dandruffy
- |
  dandy
- |
  dandyism
- |
  danger
- |
  dangerous
- |
  dangerously
- |
  dangle
- |
  dangler
- |
  dangling
- |
  Daniel
- |
  Danielle
- |
  danio
- |
  Danish
- |
  danish
- |
  dankly
- |
  dankness
- |
  Danny
- |
  danseur
- |
  danseuse
- |
  Dante
- |
  Dantean
- |
  Dantesque
- |
  Danton
- |
  Danube
- |
  Danubian
- |
  Danzig
- |
  Daphne
- |
  dapper
- |
  dapperly
- |
  dapperness
- |
  dapple
- |
  dappled
- |
  Dardanelles
- |
  daredevil
- |
  daredevilry
- |
  darer
- |
  daresay
- |
  daring
- |
  daringly
- |
  daringness
- |
  Darius
- |
  darken
- |
  darkened
- |
  darkener
- |
  darkish
- |
  darkling
- |
  darkly
- |
  darkness
- |
  darkroom
- |
  Darla
- |
  Darlene
- |
  Darling
- |
  darling
- |
  darned
- |
  darner
- |
  darning
- |
  Darold
- |
  Darrel
- |
  Darrell
- |
  Darrow
- |
  Darryl
- |
  dartboard
- |
  darter
- |
  darts
- |
  Darvon
- |
  Darwin
- |
  Darwinian
- |
  Darwinism
- |
  Darwinist
- |
  Darwinistic
- |
  Daryl
- |
  dashboard
- |
  dasher
- |
  dashiki
- |
  dashing
- |
  dashingly
- |
  dastard
- |
  dastardly
- |
  databank
- |
  database
- |
  datable
- |
  datcha
- |
  dateable
- |
  dated
- |
  datedness
- |
  dateless
- |
  dateline
- |
  dater
- |
  dative
- |
  datum
- |
  dauber
- |
  Daudet
- |
  daughter
- |
  daughterly
- |
  Daumier
- |
  daunt
- |
  daunting
- |
  dauntingly
- |
  dauntless
- |
  dauntlessly
- |
  dauphin
- |
  dauphine
- |
  Davao
- |
  Davenport
- |
  davenport
- |
  David
- |
  Davis
- |
  davit
- |
  dawdle
- |
  dawdler
- |
  Dawes
- |
  dawning
- |
  Dayan
- |
  daybed
- |
  daybook
- |
  daybreak
- |
  daycare
- |
  daydream
- |
  daydreamer
- |
  daylight
- |
  daylights
- |
  daytime
- |
  Dayton
- |
  dazed
- |
  dazedly
- |
  dazzle
- |
  dazzler
- |
  dazzling
- |
  dazzlingly
- |
  deacon
- |
  deaconate
- |
  deaconess
- |
  deaconry
- |
  deaconship
- |
  deactivate
- |
  deactivation
- |
  deadbeat
- |
  deadbolt
- |
  deaden
- |
  deadeye
- |
  Deadhead
- |
  deadhead
- |
  deadline
- |
  deadliness
- |
  deadlock
- |
  deadlocked
- |
  deadly
- |
  deadness
- |
  deadpan
- |
  deadweight
- |
  deadwood
- |
  deafen
- |
  deafening
- |
  deafeningly
- |
  deafly
- |
  deafness
- |
  dealer
- |
  dealership
- |
  dealing
- |
  dealings
- |
  dealt
- |
  Deane
- |
  deanery
- |
  Deanna
- |
  Deanne
- |
  deanship
- |
  Dearborn
- |
  dearest
- |
  dearly
- |
  dearness
- |
  dearth
- |
  death
- |
  deathbed
- |
  deathblow
- |
  deathless
- |
  deathlessly
- |
  deathlike
- |
  deathly
- |
  deathtrap
- |
  deathwatch
- |
  debacle
- |
  debar
- |
  debark
- |
  debarkation
- |
  debarment
- |
  debase
- |
  debasement
- |
  debaser
- |
  debatable
- |
  debate
- |
  debater
- |
  debating
- |
  debauch
- |
  debauched
- |
  debauchee
- |
  debaucher
- |
  debauchery
- |
  Debbie
- |
  Debby
- |
  debenture
- |
  debilitate
- |
  debilitated
- |
  debilitating
- |
  debilitation
- |
  debilitative
- |
  debility
- |
  debit
- |
  debonair
- |
  debonaire
- |
  debonairly
- |
  Debora
- |
  Deborah
- |
  debouch
- |
  debouchment
- |
  Debra
- |
  Debrecen
- |
  debridement
- |
  debrief
- |
  debriefing
- |
  debris
- |
  debtor
- |
  debug
- |
  debugger
- |
  debunk
- |
  debunker
- |
  Debussy
- |
  debut
- |
  debutante
- |
  decade
- |
  decadence
- |
  decadent
- |
  decadently
- |
  decaf
- |
  decaffeinate
- |
  decagon
- |
  decagonal
- |
  decagonally
- |
  decagram
- |
  decahedra
- |
  decahedral
- |
  decahedron
- |
  decal
- |
  decalcifier
- |
  decalcify
- |
  decalcomania
- |
  decaliter
- |
  Decalog
- |
  Decalogue
- |
  decameter
- |
  decamp
- |
  decampment
- |
  decant
- |
  decantation
- |
  decanter
- |
  decapitate
- |
  decapitation
- |
  decapitator
- |
  decasyllabic
- |
  decasyllable
- |
  decathlete
- |
  decathlon
- |
  Decatur
- |
  decay
- |
  decayed
- |
  Deccan
- |
  decease
- |
  deceased
- |
  decedent
- |
  deceit
- |
  deceitful
- |
  deceitfully
- |
  deceive
- |
  deceiver
- |
  deceivingly
- |
  decelerate
- |
  deceleration
- |
  decelerator
- |
  December
- |
  decency
- |
  decennial
- |
  decennially
- |
  decent
- |
  decently
- |
  decentness
- |
  decentralize
- |
  deception
- |
  deceptive
- |
  deceptively
- |
  decibel
- |
  decidable
- |
  decide
- |
  decided
- |
  decidedly
- |
  decidedness
- |
  decider
- |
  deciduous
- |
  deciduously
- |
  decigram
- |
  deciliter
- |
  decillion
- |
  decillionth
- |
  decimal
- |
  decimally
- |
  decimate
- |
  decimation
- |
  decimator
- |
  decimeter
- |
  decipher
- |
  decipherable
- |
  decipherment
- |
  decision
- |
  decisive
- |
  decisively
- |
  decisiveness
- |
  deckhand
- |
  declaim
- |
  declaimer
- |
  declamation
- |
  declamatory
- |
  declaration
- |
  declarative
- |
  declaratory
- |
  declare
- |
  declarer
- |
  declasse
- |
  declassee
- |
  declassify
- |
  declension
- |
  declensional
- |
  declinable
- |
  declination
- |
  decline
- |
  decliner
- |
  declivitous
- |
  declivity
- |
  decoct
- |
  decoction
- |
  decode
- |
  decoder
- |
  decolletage
- |
  decollete
- |
  decolletee
- |
  decolonize
- |
  decommission
- |
  decomposable
- |
  decompose
- |
  decomposed
- |
  decomposer
- |
  decompress
- |
  decongest
- |
  decongestant
- |
  decongestion
- |
  decongestive
- |
  deconstruct
- |
  decontrol
- |
  decor
- |
  decorate
- |
  decorating
- |
  decoration
- |
  decorative
- |
  decoratively
- |
  decorator
- |
  decorous
- |
  decorously
- |
  decorousness
- |
  decorum
- |
  decorums
- |
  decoupage
- |
  decoy
- |
  decoyer
- |
  decrease
- |
  decreasingly
- |
  decree
- |
  decrement
- |
  decremental
- |
  decrepit
- |
  decrepitly
- |
  decrepitude
- |
  decrescendo
- |
  decretal
- |
  decrier
- |
  decry
- |
  decussate
- |
  decussation
- |
  dedicate
- |
  dedicated
- |
  dedication
- |
  dedicative
- |
  dedicator
- |
  dedicatory
- |
  deduce
- |
  deducible
- |
  deduct
- |
  deductible
- |
  deduction
- |
  deductive
- |
  deductively
- |
  deejay
- |
  Deena
- |
  deepen
- |
  deepfreeze
- |
  deepfroze
- |
  deepfrozen
- |
  deeply
- |
  deepness
- |
  deerfly
- |
  deerskin
- |
  deescalate
- |
  deescalation
- |
  deface
- |
  defacement
- |
  defacer
- |
  defalcate
- |
  defalcation
- |
  defalcator
- |
  defamation
- |
  defamatory
- |
  defame
- |
  defamer
- |
  default
- |
  defaulter
- |
  defeasance
- |
  defeat
- |
  defeater
- |
  defeatism
- |
  defeatist
- |
  defecate
- |
  defecation
- |
  defecator
- |
  defecatory
- |
  defect
- |
  defection
- |
  defective
- |
  defectively
- |
  defector
- |
  defence
- |
  defend
- |
  defendable
- |
  defendant
- |
  defender
- |
  defenestrate
- |
  defense
- |
  defenseless
- |
  defensible
- |
  defensibly
- |
  defensive
- |
  defensively
- |
  defer
- |
  deference
- |
  deferential
- |
  deferment
- |
  deferrable
- |
  deferral
- |
  deferrer
- |
  defiance
- |
  defiant
- |
  defiantly
- |
  defibrillate
- |
  deficiency
- |
  deficient
- |
  deficiently
- |
  deficit
- |
  defier
- |
  defile
- |
  defilement
- |
  defiler
- |
  definable
- |
  definably
- |
  define
- |
  defined
- |
  definer
- |
  definite
- |
  definitely
- |
  definiteness
- |
  definition
- |
  definitive
- |
  definitively
- |
  deflagrate
- |
  deflagration
- |
  deflagrator
- |
  deflate
- |
  deflated
- |
  deflation
- |
  deflationary
- |
  deflationist
- |
  deflator
- |
  deflect
- |
  deflectable
- |
  deflection
- |
  deflective
- |
  deflector
- |
  defloration
- |
  deflower
- |
  deflowered
- |
  Defoe
- |
  defog
- |
  defogger
- |
  defoliant
- |
  defoliate
- |
  defoliation
- |
  defoliator
- |
  deforest
- |
  deform
- |
  deformable
- |
  deformation
- |
  deformed
- |
  deformity
- |
  defraud
- |
  defraudation
- |
  defrauder
- |
  defray
- |
  defrayable
- |
  defrayal
- |
  defrayment
- |
  defrock
- |
  defrost
- |
  defroster
- |
  deftly
- |
  deftness
- |
  defunct
- |
  defuse
- |
  degage
- |
  Degas
- |
  degas
- |
  degauss
- |
  degausser
- |
  degaussing
- |
  degeneracy
- |
  degenerate
- |
  degenerately
- |
  degeneration
- |
  degenerative
- |
  degradable
- |
  degradation
- |
  degradative
- |
  degrade
- |
  degraded
- |
  degrader
- |
  degrading
- |
  degree
- |
  dehisce
- |
  dehiscence
- |
  dehiscent
- |
  dehorn
- |
  dehumanize
- |
  dehumidifier
- |
  dehumidify
- |
  dehydrate
- |
  dehydrated
- |
  dehydration
- |
  dehydrator
- |
  deice
- |
  deicer
- |
  deification
- |
  deify
- |
  deign
- |
  deionize
- |
  Deirdre
- |
  deism
- |
  deist
- |
  deistic
- |
  deistical
- |
  deistically
- |
  Deity
- |
  deity
- |
  deject
- |
  dejected
- |
  dejectedly
- |
  dejectedness
- |
  dejection
- |
  dekagram
- |
  dekaliter
- |
  dekameter
- |
  Delacroix
- |
  Delano
- |
  Delaware
- |
  Delawarean
- |
  Delawarian
- |
  delay
- |
  delayed
- |
  delayer
- |
  Delbert
- |
  delectable
- |
  delectably
- |
  delectation
- |
  delegable
- |
  delegate
- |
  delegation
- |
  delegator
- |
  delete
- |
  deleterious
- |
  deletion
- |
  delft
- |
  delftware
- |
  Delhi
- |
  Delia
- |
  Delian
- |
  deliberate
- |
  deliberately
- |
  deliberation
- |
  deliberative
- |
  deliberator
- |
  Delibes
- |
  delicacy
- |
  delicate
- |
  delicately
- |
  delicateness
- |
  delicatessen
- |
  delicious
- |
  deliciously
- |
  delict
- |
  delight
- |
  delighted
- |
  delightedly
- |
  delightful
- |
  delightfully
- |
  Delilah
- |
  delimit
- |
  delimitation
- |
  delimiter
- |
  delineate
- |
  delineation
- |
  delineative
- |
  delineator
- |
  delinquency
- |
  delinquent
- |
  delinquently
- |
  deliquesce
- |
  deliquescent
- |
  deliria
- |
  delirious
- |
  deliriously
- |
  delirium
- |
  Delius
- |
  deliver
- |
  deliverable
- |
  deliverance
- |
  deliverer
- |
  delivery
- |
  deliveryman
- |
  Della
- |
  Delmar
- |
  Delmer
- |
  Delores
- |
  Delos
- |
  delouse
- |
  Delphi
- |
  delphinia
- |
  delphinium
- |
  Delphinus
- |
  delta
- |
  deltaic
- |
  deltoid
- |
  delude
- |
  deluded
- |
  deludedly
- |
  deluder
- |
  Deluge
- |
  deluge
- |
  delusion
- |
  delusional
- |
  delusive
- |
  delusively
- |
  delusiveness
- |
  deluxe
- |
  delve
- |
  delver
- |
  demagnetize
- |
  demagnetizer
- |
  demagog
- |
  demagogic
- |
  demagogical
- |
  demagogue
- |
  demagoguery
- |
  demagogy
- |
  demand
- |
  demandable
- |
  demander
- |
  demanding
- |
  demandingly
- |
  demands
- |
  demarcate
- |
  demarcation
- |
  demarcative
- |
  demarcator
- |
  demarche
- |
  demean
- |
  demeaning
- |
  demeanor
- |
  demeanour
- |
  demented
- |
  dementedly
- |
  dementia
- |
  demerit
- |
  Demerol
- |
  demesne
- |
  Demeter
- |
  demigod
- |
  demigoddess
- |
  demijohn
- |
  demilitarize
- |
  demimondaine
- |
  demimonde
- |
  demineralize
- |
  demise
- |
  demission
- |
  demit
- |
  demitasse
- |
  demiurge
- |
  demiurgic
- |
  demiurgical
- |
  demobilise
- |
  demobilize
- |
  democracy
- |
  Democrat
- |
  democrat
- |
  Democratic
- |
  democratic
- |
  democratize
- |
  Democritus
- |
  demode
- |
  demodulate
- |
  demodulation
- |
  demodulator
- |
  demographer
- |
  demographic
- |
  demographics
- |
  demography
- |
  demoiselle
- |
  demolish
- |
  demolition
- |
  demon
- |
  demonetize
- |
  demoniac
- |
  demoniacal
- |
  demoniacally
- |
  demonic
- |
  demonical
- |
  demonically
- |
  demonization
- |
  demonize
- |
  demonologist
- |
  demonology
- |
  demonstrable
- |
  demonstrably
- |
  demonstrate
- |
  demonstrator
- |
  demoralize
- |
  demoralized
- |
  demoralizer
- |
  demoralizing
- |
  Demosthenes
- |
  demote
- |
  Demotic
- |
  demotic
- |
  demotion
- |
  Dempsey
- |
  demulcent
- |
  demur
- |
  demure
- |
  demurely
- |
  demureness
- |
  demurral
- |
  demurrer
- |
  demystify
- |
  Denali
- |
  denar
- |
  denari
- |
  denaturant
- |
  denaturation
- |
  denature
- |
  denatured
- |
  dendrite
- |
  dendrologist
- |
  dendrology
- |
  Deneb
- |
  Denebola
- |
  dengue
- |
  deniability
- |
  deniable
- |
  deniably
- |
  denial
- |
  denier
- |
  denigrate
- |
  denigration
- |
  denigrator
- |
  denigratory
- |
  denim
- |
  denims
- |
  Denis
- |
  Denise
- |
  denizen
- |
  denizenship
- |
  Denmark
- |
  Dennis
- |
  Denny
- |
  denominate
- |
  denomination
- |
  denominator
- |
  denotation
- |
  denotational
- |
  denotative
- |
  denotatively
- |
  denote
- |
  denouement
- |
  denounce
- |
  denouncement
- |
  denouncer
- |
  Denpasar
- |
  dense
- |
  densely
- |
  denseness
- |
  density
- |
  dental
- |
  dentally
- |
  dentate
- |
  dented
- |
  dentifrice
- |
  dentin
- |
  dentinal
- |
  dentine
- |
  dentist
- |
  dentistry
- |
  dentition
- |
  Denton
- |
  denture
- |
  dentures
- |
  denuclearize
- |
  denudation
- |
  denude
- |
  denunciation
- |
  denunciative
- |
  denunciatory
- |
  Denver
- |
  deodar
- |
  deodorant
- |
  deodorize
- |
  deodorizer
- |
  deoxidize
- |
  deoxyribose
- |
  depart
- |
  departed
- |
  departee
- |
  department
- |
  departmental
- |
  departure
- |
  depend
- |
  dependable
- |
  dependably
- |
  dependance
- |
  dependancy
- |
  dependant
- |
  dependence
- |
  dependency
- |
  dependent
- |
  dependently
- |
  depict
- |
  depicter
- |
  depiction
- |
  depictor
- |
  depilatory
- |
  deplane
- |
  deplete
- |
  depleted
- |
  depletion
- |
  deplorable
- |
  deplorably
- |
  deplore
- |
  deploring
- |
  deploy
- |
  deployable
- |
  deployment
- |
  depolarize
- |
  depoliticize
- |
  deponent
- |
  depopulate
- |
  depopulation
- |
  deport
- |
  deportable
- |
  deportation
- |
  deportee
- |
  deportment
- |
  depose
- |
  deposit
- |
  deposition
- |
  depositional
- |
  depositor
- |
  depository
- |
  depot
- |
  deprave
- |
  depraved
- |
  depravity
- |
  deprecate
- |
  deprecating
- |
  deprecation
- |
  deprecative
- |
  deprecator
- |
  deprecatory
- |
  depreciate
- |
  depreciation
- |
  depreciative
- |
  depreciator
- |
  depreciatory
- |
  depredate
- |
  depredation
- |
  depredations
- |
  depredator
- |
  depredatory
- |
  depress
- |
  depressant
- |
  depressed
- |
  depressing
- |
  depressingly
- |
  depression
- |
  depressive
- |
  depressively
- |
  depressor
- |
  depressurize
- |
  deprivation
- |
  deprive
- |
  deprived
- |
  deprogram
- |
  deprogrammer
- |
  depth
- |
  depths
- |
  deputation
- |
  depute
- |
  deputize
- |
  deputy
- |
  deracinate
- |
  deracinated
- |
  deracination
- |
  derail
- |
  derailleur
- |
  derailment
- |
  Derain
- |
  derange
- |
  deranged
- |
  derangement
- |
  Derby
- |
  derby
- |
  Derbyshire
- |
  deregulate
- |
  deregulation
- |
  deregulatory
- |
  Derek
- |
  derelict
- |
  dereliction
- |
  deride
- |
  derisible
- |
  derision
- |
  derisive
- |
  derisively
- |
  derisiveness
- |
  derisory
- |
  derivable
- |
  derivation
- |
  derivational
- |
  derivative
- |
  derivatively
- |
  derivatives
- |
  derive
- |
  derma
- |
  dermabrasion
- |
  dermal
- |
  dermatitis
- |
  dermatology
- |
  dermis
- |
  derogate
- |
  derogation
- |
  derogative
- |
  derogatorily
- |
  derogatory
- |
  derrick
- |
  derriere
- |
  derringer
- |
  Derry
- |
  dervish
- |
  desalinate
- |
  desalination
- |
  desalinator
- |
  desalinize
- |
  desalt
- |
  desalter
- |
  descant
- |
  Descartes
- |
  descend
- |
  descendant
- |
  descended
- |
  descendent
- |
  descent
- |
  describable
- |
  describe
- |
  describer
- |
  description
- |
  descriptive
- |
  descry
- |
  desecrate
- |
  desecrater
- |
  desecration
- |
  desecrator
- |
  desegregate
- |
  desegregated
- |
  desensitize
- |
  desensitizer
- |
  desert
- |
  deserted
- |
  deserter
- |
  desertion
- |
  deserts
- |
  deserve
- |
  deserved
- |
  deservedly
- |
  deserving
- |
  deservingly
- |
  desex
- |
  desexed
- |
  deshabille
- |
  desiccant
- |
  desiccate
- |
  desiccated
- |
  desiccation
- |
  desiccative
- |
  desiccator
- |
  desiderata
- |
  desiderative
- |
  desideratum
- |
  design
- |
  designate
- |
  designation
- |
  designative
- |
  designer
- |
  designing
- |
  designs
- |
  desirability
- |
  desirable
- |
  desirably
- |
  desire
- |
  desirer
- |
  desirous
- |
  desist
- |
  desktop
- |
  desolate
- |
  desolated
- |
  desolately
- |
  desolateness
- |
  desolating
- |
  desolation
- |
  desolator
- |
  despair
- |
  despairingly
- |
  despatch
- |
  desperado
- |
  desperate
- |
  desperately
- |
  desperation
- |
  despicable
- |
  despicably
- |
  despise
- |
  despiser
- |
  despite
- |
  despoil
- |
  despoiler
- |
  despoilment
- |
  despoliation
- |
  despond
- |
  despondence
- |
  despondency
- |
  despondent
- |
  despondently
- |
  despondingly
- |
  despot
- |
  despotic
- |
  despotically
- |
  despotism
- |
  dessert
- |
  destabilize
- |
  destination
- |
  destine
- |
  destined
- |
  destiny
- |
  destitute
- |
  destitution
- |
  destroy
- |
  destroyer
- |
  destruct
- |
  destructible
- |
  destruction
- |
  destructive
- |
  desuetude
- |
  desultorily
- |
  desultory
- |
  detach
- |
  detachable
- |
  detached
- |
  detachment
- |
  detail
- |
  detailed
- |
  detain
- |
  detainee
- |
  detainment
- |
  detect
- |
  detectable
- |
  detecter
- |
  detectible
- |
  detection
- |
  detective
- |
  detector
- |
  detente
- |
  detention
- |
  deter
- |
  detergent
- |
  deteriorate
- |
  determent
- |
  determinable
- |
  determinably
- |
  determinacy
- |
  determinant
- |
  determinate
- |
  determine
- |
  determined
- |
  determinedly
- |
  determiner
- |
  determinism
- |
  determinist
- |
  deterrence
- |
  deterrent
- |
  detest
- |
  detestable
- |
  detestably
- |
  detestation
- |
  dethrone
- |
  dethronement
- |
  detonate
- |
  detonation
- |
  detonator
- |
  detour
- |
  detox
- |
  detoxify
- |
  detract
- |
  detraction
- |
  detractive
- |
  detractor
- |
  detrain
- |
  detriment
- |
  detrimental
- |
  detrital
- |
  detritus
- |
  Detroit
- |
  detumesce
- |
  detumescence
- |
  detumescent
- |
  deuce
- |
  deuterium
- |
  Deuteronomy
- |
  deutschemark
- |
  Deutschmark
- |
  devaluate
- |
  devaluation
- |
  devalue
- |
  devalued
- |
  devastate
- |
  devastated
- |
  devastating
- |
  devastation
- |
  devastator
- |
  develop
- |
  developed
- |
  developer
- |
  developing
- |
  development
- |
  deviance
- |
  deviancy
- |
  deviant
- |
  deviate
- |
  deviation
- |
  deviationism
- |
  deviationist
- |
  deviator
- |
  device
- |
  Devil
- |
  devil
- |
  devilish
- |
  devilishly
- |
  devilishness
- |
  devilment
- |
  devilry
- |
  deviltry
- |
  devious
- |
  deviously
- |
  deviousness
- |
  devisable
- |
  devise
- |
  devisee
- |
  deviser
- |
  devisor
- |
  devitalize
- |
  devoid
- |
  devoir
- |
  devolution
- |
  devolve
- |
  devolved
- |
  devolvement
- |
  Devon
- |
  Devonian
- |
  Devonshire
- |
  devote
- |
  devoted
- |
  devotedly
- |
  devotee
- |
  devotion
- |
  devotional
- |
  devotions
- |
  devour
- |
  devourer
- |
  devout
- |
  devoutly
- |
  devoutness
- |
  dewberry
- |
  dewclaw
- |
  dewdrop
- |
  Dewey
- |
  dewily
- |
  dewiness
- |
  Dewitt
- |
  dewlap
- |
  Dexter
- |
  dexter
- |
  dexterity
- |
  dexterous
- |
  dexterously
- |
  dextral
- |
  dextrality
- |
  dextrally
- |
  dextrin
- |
  dextrose
- |
  dextrous
- |
  dextrously
- |
  dextrousness
- |
  Dhaka
- |
  dharma
- |
  Dhaulagiri
- |
  dhoti
- |
  dhurrie
- |
  diabetes
- |
  diabetic
- |
  diabolic
- |
  diabolical
- |
  diabolically
- |
  diacritic
- |
  diacritical
- |
  diadem
- |
  diademed
- |
  diaereses
- |
  diaeresis
- |
  Diaghilev
- |
  diagnose
- |
  diagnoses
- |
  diagnosis
- |
  diagnostic
- |
  diagnostics
- |
  diagonal
- |
  diagonally
- |
  diagram
- |
  diagrammable
- |
  diagrammatic
- |
  dialect
- |
  dialectal
- |
  dialectic
- |
  dialectical
- |
  dialectics
- |
  dialer
- |
  dialog
- |
  dialogue
- |
  dialyses
- |
  dialysis
- |
  dialytic
- |
  dialyze
- |
  diamagnetic
- |
  diamagnetism
- |
  diameter
- |
  diametric
- |
  diametrical
- |
  diamond
- |
  diamondback
- |
  Diana
- |
  Diane
- |
  Diann
- |
  Dianna
- |
  Dianne
- |
  dianthus
- |
  diapason
- |
  diaper
- |
  diaphanous
- |
  diaphanously
- |
  diaphoresis
- |
  diaphoretic
- |
  diaphragm
- |
  diarist
- |
  diarrhea
- |
  diarrheal
- |
  diarrheic
- |
  diarrhoea
- |
  diary
- |
  diaspora
- |
  diastase
- |
  diastole
- |
  diastolic
- |
  diathermic
- |
  diathermy
- |
  diatom
- |
  diatomaceous
- |
  diatomic
- |
  diatonic
- |
  diatonically
- |
  diatonicism
- |
  diatribe
- |
  diazepam
- |
  dibble
- |
  dicer
- |
  dicey
- |
  dichotomize
- |
  dichotomous
- |
  dichotomy
- |
  Dickens
- |
  Dickensian
- |
  dicker
- |
  dickey
- |
  dickie
- |
  Dickinson
- |
  dicky
- |
  dicot
- |
  dicotyledon
- |
  dicta
- |
  Dictaphone
- |
  dictate
- |
  dictation
- |
  dictator
- |
  dictatorial
- |
  dictatorship
- |
  diction
- |
  dictionary
- |
  dictum
- |
  didactic
- |
  didactical
- |
  didactically
- |
  didacticism
- |
  diddle
- |
  diddler
- |
  Diderot
- |
  Didrikson
- |
  didst
- |
  Diefenbaker
- |
  diehard
- |
  dielectric
- |
  Dienbienphu
- |
  diereses
- |
  dieresis
- |
  diesel
- |
  dieseling
- |
  dieselize
- |
  dietary
- |
  dieter
- |
  dietetic
- |
  dietetics
- |
  dietician
- |
  dieting
- |
  dietitian
- |
  Dietrich
- |
  differ
- |
  difference
- |
  different
- |
  differential
- |
  differently
- |
  difficult
- |
  difficulties
- |
  difficultly
- |
  difficulty
- |
  diffidence
- |
  diffident
- |
  diffidently
- |
  diffract
- |
  diffraction
- |
  diffractive
- |
  diffuse
- |
  diffusely
- |
  diffuseness
- |
  diffusible
- |
  diffusion
- |
  diffusive
- |
  digerati
- |
  digest
- |
  digestible
- |
  digestion
- |
  digestive
- |
  digger
- |
  digit
- |
  digital
- |
  digitalis
- |
  digitally
- |
  digitigrade
- |
  digitization
- |
  digitize
- |
  dignified
- |
  dignify
- |
  dignitary
- |
  dignity
- |
  digraph
- |
  digraphic
- |
  digress
- |
  digresser
- |
  digression
- |
  digressive
- |
  digressively
- |
  Dijon
- |
  dilapidated
- |
  dilapidation
- |
  dilatable
- |
  dilatation
- |
  dilate
- |
  dilated
- |
  dilation
- |
  dilator
- |
  dilatorily
- |
  dilatoriness
- |
  dilatory
- |
  dilemma
- |
  dilettante
- |
  dilettanti
- |
  dilettantish
- |
  dilettantism
- |
  diligence
- |
  diligent
- |
  diligently
- |
  Dillinger
- |
  dilly
- |
  dillydally
- |
  diluent
- |
  dilute
- |
  diluter
- |
  dilution
- |
  DiMaggio
- |
  dimension
- |
  dimensional
- |
  dimensions
- |
  diminish
- |
  diminishable
- |
  diminishment
- |
  diminuendi
- |
  diminuendo
- |
  diminution
- |
  diminutive
- |
  diminutively
- |
  dimity
- |
  dimly
- |
  dimmer
- |
  dimness
- |
  dimorphic
- |
  dimorphism
- |
  dimple
- |
  dimpled
- |
  dimply
- |
  dimwit
- |
  dimwitted
- |
  Dinah
- |
  dinar
- |
  diner
- |
  Dinesen
- |
  dinette
- |
  dinghy
- |
  dingily
- |
  dinginess
- |
  dingle
- |
  dingo
- |
  dingus
- |
  dingy
- |
  dinky
- |
  dinner
- |
  dinnertime
- |
  dinnerware
- |
  dinosaur
- |
  diocesan
- |
  diocese
- |
  Diocletian
- |
  diode
- |
  Diogenes
- |
  Dionysiac
- |
  Dionysian
- |
  dionysian
- |
  Dionysius
- |
  Dionysos
- |
  Dionysus
- |
  diorama
- |
  dioxide
- |
  dioxin
- |
  diphtheria
- |
  diphtherial
- |
  diphtheric
- |
  diphtheritic
- |
  diphthong
- |
  diphthongal
- |
  diploid
- |
  diploma
- |
  diplomacy
- |
  diplomat
- |
  diplomatic
- |
  diplomatist
- |
  dipolar
- |
  dipole
- |
  dipper
- |
  dipping
- |
  dipsomania
- |
  dipsomaniac
- |
  dipstick
- |
  dipteran
- |
  dipterous
- |
  diptych
- |
  direct
- |
  direction
- |
  directional
- |
  directions
- |
  directive
- |
  directly
- |
  directness
- |
  director
- |
  directorate
- |
  directorial
- |
  directorship
- |
  directory
- |
  direful
- |
  direfully
- |
  direly
- |
  direness
- |
  dirge
- |
  dirgeful
- |
  dirham
- |
  dirigible
- |
  dirndl
- |
  dirtily
- |
  dirtiness
- |
  dirty
- |
  disability
- |
  disable
- |
  disabled
- |
  disablement
- |
  disabling
- |
  disabuse
- |
  disaccharide
- |
  disadvantage
- |
  disaffect
- |
  disaffected
- |
  disaffection
- |
  disaffiliate
- |
  disagree
- |
  disagreeable
- |
  disagreeably
- |
  disagreement
- |
  disallow
- |
  disallowance
- |
  disappear
- |
  disappoint
- |
  disappointed
- |
  disapproval
- |
  disapprove
- |
  disarm
- |
  disarmament
- |
  disarming
- |
  disarmingly
- |
  disarrange
- |
  disarray
- |
  disassemble
- |
  disassociate
- |
  disaster
- |
  disastrous
- |
  disastrously
- |
  disavow
- |
  disavowal
- |
  disband
- |
  disbandment
- |
  disbar
- |
  disbarment
- |
  disbelief
- |
  disbelieve
- |
  disbeliever
- |
  disbelieving
- |
  disburden
- |
  disbursal
- |
  disburse
- |
  disbursement
- |
  disburser
- |
  discard
- |
  discern
- |
  discerner
- |
  discernible
- |
  discernibly
- |
  discerning
- |
  discerningly
- |
  discernment
- |
  discharge
- |
  Disciple
- |
  disciple
- |
  discipleship
- |
  disciplinary
- |
  discipline
- |
  disciplined
- |
  disclaim
- |
  disclaimer
- |
  disclose
- |
  discloser
- |
  disclosure
- |
  disco
- |
  discolor
- |
  discolour
- |
  discomfit
- |
  discomfiture
- |
  discomfort
- |
  discommode
- |
  discompose
- |
  discomposure
- |
  disconcert
- |
  disconcerted
- |
  disconnect
- |
  disconnected
- |
  disconsolate
- |
  discontent
- |
  discontented
- |
  discontinue
- |
  discord
- |
  discordance
- |
  discordant
- |
  discordantly
- |
  discotheque
- |
  discount
- |
  discountable
- |
  discounted
- |
  discounter
- |
  discourage
- |
  discouraged
- |
  discouraging
- |
  discourse
- |
  discourteous
- |
  discourtesy
- |
  discover
- |
  discoverable
- |
  discoverer
- |
  discovery
- |
  discredit
- |
  discredited
- |
  discreet
- |
  discreetly
- |
  discreetness
- |
  discrepancy
- |
  discrepant
- |
  discrete
- |
  discretely
- |
  discreteness
- |
  discretion
- |
  discriminant
- |
  discriminate
- |
  discursive
- |
  discursively
- |
  discus
- |
  discuss
- |
  discussant
- |
  discussion
- |
  disdain
- |
  disdainful
- |
  disdainfully
- |
  disease
- |
  diseased
- |
  disembark
- |
  disembodied
- |
  disembody
- |
  disembogue
- |
  disembowel
- |
  disenchant
- |
  disenchanted
- |
  disencumber
- |
  disengage
- |
  disentangle
- |
  disentangler
- |
  disestablish
- |
  disesteem
- |
  disfavor
- |
  disfavour
- |
  disfigure
- |
  disfigured
- |
  disfiguring
- |
  disfranchise
- |
  disgorge
- |
  disgorgement
- |
  disgrace
- |
  disgraced
- |
  disgraceful
- |
  disgruntle
- |
  disgruntled
- |
  disguise
- |
  disguised
- |
  disgust
- |
  disgusted
- |
  disgustedly
- |
  disgustful
- |
  disgusting
- |
  disgustingly
- |
  dishabille
- |
  disharmony
- |
  dishcloth
- |
  dishearten
- |
  disheartened
- |
  dished
- |
  dishes
- |
  dishevel
- |
  disheveled
- |
  dishevelled
- |
  dishevelment
- |
  dishonest
- |
  dishonestly
- |
  dishonesty
- |
  dishonor
- |
  dishonorable
- |
  dishonorably
- |
  dishpan
- |
  dishrag
- |
  dishtowel
- |
  dishwasher
- |
  dishwater
- |
  disillusion
- |
  disincline
- |
  disinclined
- |
  disinfect
- |
  disinfectant
- |
  disinfection
- |
  disinflation
- |
  disingenuity
- |
  disingenuous
- |
  disinherit
- |
  disintegrate
- |
  disinter
- |
  disinterest
- |
  disinterment
- |
  disjoin
- |
  disjoint
- |
  disjointed
- |
  disjointedly
- |
  disjunct
- |
  disjunction
- |
  disjunctive
- |
  diskette
- |
  dislike
- |
  dislocate
- |
  dislocation
- |
  dislodge
- |
  dislodgement
- |
  dislodgment
- |
  disloyal
- |
  disloyally
- |
  disloyalty
- |
  dismal
- |
  dismally
- |
  dismantle
- |
  dismantler
- |
  dismay
- |
  dismayed
- |
  dismayingly
- |
  dismember
- |
  dismiss
- |
  dismissal
- |
  dismissible
- |
  dismissive
- |
  dismissively
- |
  dismount
- |
  dismountable
- |
  Disney
- |
  disobedience
- |
  disobedient
- |
  disobey
- |
  disoblige
- |
  disorder
- |
  disordered
- |
  disorderly
- |
  disorganised
- |
  disorganize
- |
  disorganized
- |
  disorient
- |
  disoriented
- |
  disorienting
- |
  disown
- |
  disparage
- |
  disparaging
- |
  disparate
- |
  disparately
- |
  disparity
- |
  dispassion
- |
  dispatch
- |
  dispatcher
- |
  dispel
- |
  dispeller
- |
  dispensable
- |
  dispensary
- |
  dispensation
- |
  dispense
- |
  dispenser
- |
  dispersal
- |
  disperse
- |
  dispersed
- |
  disperser
- |
  dispersible
- |
  dispersion
- |
  dispersive
- |
  dispirit
- |
  dispirited
- |
  dispiritedly
- |
  dispiriting
- |
  displace
- |
  displacement
- |
  display
- |
  displease
- |
  displeased
- |
  displeasure
- |
  disport
- |
  disposable
- |
  disposal
- |
  dispose
- |
  disposed
- |
  disposer
- |
  disposition
- |
  dispossess
- |
  dispraise
- |
  dispraiser
- |
  disproof
- |
  disprovable
- |
  disproval
- |
  disprove
- |
  disputable
- |
  disputably
- |
  disputant
- |
  disputation
- |
  disputatious
- |
  dispute
- |
  disputer
- |
  disqualify
- |
  disquiet
- |
  disquieted
- |
  disquieting
- |
  disquietude
- |
  disquisition
- |
  Disraeli
- |
  disregard
- |
  disregardful
- |
  disrepair
- |
  disreputable
- |
  disreputably
- |
  disrepute
- |
  disrespect
- |
  disrobe
- |
  disrupt
- |
  disrupter
- |
  disruption
- |
  disruptive
- |
  disruptively
- |
  disruptor
- |
  dissatisfied
- |
  dissatisfy
- |
  dissect
- |
  dissected
- |
  dissection
- |
  dissector
- |
  dissemblance
- |
  dissemble
- |
  dissembler
- |
  disseminate
- |
  disseminated
- |
  disseminator
- |
  dissension
- |
  Dissent
- |
  dissent
- |
  dissenter
- |
  dissenting
- |
  dissertation
- |
  disservice
- |
  dissever
- |
  dissidence
- |
  dissident
- |
  dissimilar
- |
  dissimilarly
- |
  dissimulate
- |
  dissimulator
- |
  dissipate
- |
  dissipated
- |
  dissipater
- |
  dissipation
- |
  dissipative
- |
  dissipator
- |
  dissociate
- |
  dissociation
- |
  dissociative
- |
  dissolute
- |
  dissolutely
- |
  dissolution
- |
  dissolvable
- |
  dissolve
- |
  dissolver
- |
  dissonance
- |
  dissonant
- |
  dissonantly
- |
  dissuade
- |
  dissuader
- |
  dissuasion
- |
  dissuasive
- |
  distaff
- |
  distal
- |
  distally
- |
  distance
- |
  distanced
- |
  distant
- |
  distantly
- |
  distantness
- |
  distaste
- |
  distasteful
- |
  distemper
- |
  distempered
- |
  distend
- |
  distended
- |
  distensible
- |
  distension
- |
  distention
- |
  distich
- |
  distil
- |
  distill
- |
  distillate
- |
  distillation
- |
  distiller
- |
  distillery
- |
  distinct
- |
  distinction
- |
  distinctive
- |
  distinctly
- |
  distinctness
- |
  distingue
- |
  distinguee
- |
  distinguish
- |
  distort
- |
  distorted
- |
  distortedly
- |
  distortion
- |
  distortional
- |
  distract
- |
  distracted
- |
  distractedly
- |
  distracting
- |
  distraction
- |
  distrain
- |
  distrainer
- |
  distrainment
- |
  distrait
- |
  distraite
- |
  distraught
- |
  distress
- |
  distressed
- |
  distressful
- |
  distressing
- |
  distributary
- |
  distribute
- |
  distributed
- |
  distribution
- |
  distributive
- |
  distributor
- |
  district
- |
  distrust
- |
  distrustful
- |
  disturb
- |
  disturbance
- |
  disturbed
- |
  disturber
- |
  disturbing
- |
  disturbingly
- |
  disunite
- |
  disunity
- |
  disuse
- |
  disused
- |
  ditch
- |
  dither
- |
  dithered
- |
  ditherer
- |
  dithery
- |
  dithyramb
- |
  dithyrambic
- |
  ditsy
- |
  ditto
- |
  ditty
- |
  ditzy
- |
  diuretic
- |
  diurnal
- |
  diurnally
- |
  divagate
- |
  divagation
- |
  divalence
- |
  divalent
- |
  divan
- |
  divaricate
- |
  divarication
- |
  diver
- |
  diverge
- |
  divergence
- |
  divergency
- |
  divergent
- |
  divergently
- |
  divers
- |
  diverse
- |
  diversely
- |
  diverseness
- |
  diversify
- |
  diversion
- |
  diversionary
- |
  diversity
- |
  divert
- |
  diverter
- |
  diverticula
- |
  diverticulum
- |
  divertimenti
- |
  divertimento
- |
  diverting
- |
  divertingly
- |
  divest
- |
  divestiture
- |
  divestment
- |
  dividable
- |
  divide
- |
  dividend
- |
  dividends
- |
  divider
- |
  divination
- |
  divinatory
- |
  divine
- |
  divinely
- |
  divineness
- |
  diviner
- |
  diving
- |
  Divinity
- |
  divinity
- |
  divisibility
- |
  divisible
- |
  division
- |
  divisional
- |
  divisive
- |
  divisively
- |
  divisiveness
- |
  divisor
- |
  divorce
- |
  divorced
- |
  divorcee
- |
  divorcement
- |
  divot
- |
  divulgation
- |
  divulge
- |
  divulgence
- |
  divvy
- |
  Dixie
- |
  Dixieland
- |
  Diyarbakir
- |
  dizygotic
- |
  dizzily
- |
  dizziness
- |
  dizzy
- |
  dizzying
- |
  Djakarta
- |
  djellaba
- |
  djellabah
- |
  Djibouti
- |
  djinn
- |
  Dnepr
- |
  Dnieper
- |
  Dniester
- |
  doable
- |
  dobbin
- |
  doberman
- |
  dobra
- |
  docent
- |
  Docetism
- |
  Docetist
- |
  docile
- |
  docilely
- |
  docility
- |
  dockage
- |
  docket
- |
  dockhand
- |
  dockland
- |
  docks
- |
  dockworker
- |
  dockyard
- |
  doctor
- |
  doctoral
- |
  doctorate
- |
  doctoring
- |
  doctrinaire
- |
  doctrinal
- |
  doctrinally
- |
  doctrine
- |
  docudrama
- |
  document
- |
  documentable
- |
  documental
- |
  documentary
- |
  documenter
- |
  dodder
- |
  doddering
- |
  dodecagon
- |
  dodecahedra
- |
  dodecahedron
- |
  Dodecanese
- |
  dodge
- |
  dodger
- |
  Dodgson
- |
  dodgy
- |
  Dodoma
- |
  doeskin
- |
  dogbane
- |
  dogcart
- |
  dogcatcher
- |
  dogear
- |
  dogeared
- |
  dogfight
- |
  dogfish
- |
  dogged
- |
  doggedly
- |
  doggedness
- |
  doggerel
- |
  doggie
- |
  doggone
- |
  doggy
- |
  doghouse
- |
  dogie
- |
  dogleg
- |
  dogma
- |
  dogmata
- |
  dogmatic
- |
  dogmatically
- |
  dogmatism
- |
  dogmatist
- |
  dogtrot
- |
  dogwood
- |
  doily
- |
  doing
- |
  doings
- |
  Dolby
- |
  doldrums
- |
  doleful
- |
  dolefully
- |
  dolefulness
- |
  dollar
- |
  Dollfuss
- |
  dollish
- |
  dollop
- |
  Dolly
- |
  dolly
- |
  dolmen
- |
  dolomite
- |
  dolomitic
- |
  dolor
- |
  Dolores
- |
  dolorous
- |
  dolorously
- |
  dolorousness
- |
  dolour
- |
  dolphin
- |
  doltish
- |
  doltishness
- |
  domain
- |
  domaine
- |
  domainial
- |
  domed
- |
  domestic
- |
  domesticable
- |
  domestically
- |
  domesticate
- |
  domesticated
- |
  domesticity
- |
  domicil
- |
  domicile
- |
  domiciled
- |
  domiciliary
- |
  dominance
- |
  dominant
- |
  dominantly
- |
  dominate
- |
  domination
- |
  dominator
- |
  dominatrices
- |
  dominatrix
- |
  domineer
- |
  domineering
- |
  Domingo
- |
  Dominic
- |
  Dominica
- |
  Dominican
- |
  Dominick
- |
  dominie
- |
  Dominion
- |
  dominion
- |
  dominions
- |
  Domino
- |
  domino
- |
  dominoes
- |
  dominos
- |
  Domitian
- |
  Donal
- |
  Donald
- |
  donate
- |
  Donatello
- |
  donation
- |
  donative
- |
  donator
- |
  Donbas
- |
  Donetsk
- |
  dongle
- |
  Donizetti
- |
  donjon
- |
  donkey
- |
  Donna
- |
  Donne
- |
  donne
- |
  donnee
- |
  Donnie
- |
  donnybrook
- |
  donor
- |
  Donovan
- |
  donut
- |
  doodad
- |
  doodle
- |
  doodlebug
- |
  doodler
- |
  doohickey
- |
  doomed
- |
  doomsayer
- |
  doomsday
- |
  doorbell
- |
  doorjamb
- |
  doorkeeper
- |
  doorknob
- |
  doorman
- |
  doormat
- |
  doorplate
- |
  doorstep
- |
  doorstop
- |
  doorway
- |
  dooryard
- |
  doozie
- |
  doozy
- |
  dopamine
- |
  doper
- |
  dopester
- |
  dopey
- |
  dopily
- |
  dopiness
- |
  doping
- |
  doppelganger
- |
  Dorado
- |
  Dorchester
- |
  Doreen
- |
  Doric
- |
  Doris
- |
  dorky
- |
  dormancy
- |
  dormant
- |
  dormer
- |
  dormice
- |
  dormitory
- |
  dormouse
- |
  Dorothea
- |
  Dorothy
- |
  dorsal
- |
  dorsally
- |
  Dorset
- |
  Dorsetshire
- |
  Dortmund
- |
  dosage
- |
  dosimeter
- |
  dosimetry
- |
  dossier
- |
  Dostoevski
- |
  Dostoevsky
- |
  Dostoyevski
- |
  Dostoyevsky
- |
  dotage
- |
  dotard
- |
  doter
- |
  doting
- |
  dotingly
- |
  dotted
- |
  dotter
- |
  Dottie
- |
  Dotty
- |
  dotty
- |
  Douala
- |
  double
- |
  doubleheader
- |
  doubles
- |
  doublespeak
- |
  doublet
- |
  doublethink
- |
  doublets
- |
  doubloon
- |
  doubly
- |
  doubt
- |
  doubtable
- |
  doubter
- |
  doubtful
- |
  doubtfully
- |
  doubtfulness
- |
  doubtingly
- |
  doubtless
- |
  doubtlessly
- |
  douche
- |
  dough
- |
  doughboy
- |
  doughiness
- |
  doughnut
- |
  doughty
- |
  doughy
- |
  Douglas
- |
  Douglass
- |
  dourly
- |
  dourness
- |
  Douro
- |
  douse
- |
  douser
- |
  dovecote
- |
  Dover
- |
  dovetail
- |
  dovish
- |
  dovishness
- |
  dowager
- |
  dowdily
- |
  dowdiness
- |
  dowdy
- |
  dowel
- |
  dower
- |
  dowitcher
- |
  downbeat
- |
  downburst
- |
  downcast
- |
  downdraft
- |
  downer
- |
  downfall
- |
  downfallen
- |
  downgrade
- |
  downhearted
- |
  downhill
- |
  downing
- |
  download
- |
  downloadable
- |
  Downpatrick
- |
  downplay
- |
  downpour
- |
  downrange
- |
  downright
- |
  downriver
- |
  downs
- |
  downscale
- |
  downshift
- |
  downside
- |
  downsize
- |
  downsizing
- |
  downspout
- |
  downstage
- |
  downstairs
- |
  downstate
- |
  downstream
- |
  downstroke
- |
  downswing
- |
  downtick
- |
  downtime
- |
  downtown
- |
  downtrodden
- |
  downturn
- |
  downward
- |
  downwardly
- |
  downwards
- |
  downwind
- |
  downy
- |
  dowry
- |
  dowse
- |
  dowser
- |
  dowsing
- |
  doxological
- |
  doxology
- |
  doyen
- |
  doyenne
- |
  Doyle
- |
  doyley
- |
  dozen
- |
  dozens
- |
  dozenth
- |
  dozer
- |
  drably
- |
  drabness
- |
  drachma
- |
  drachmae
- |
  drachmai
- |
  Draco
- |
  Draconian
- |
  draconian
- |
  draconic
- |
  Dracula
- |
  draft
- |
  draftee
- |
  drafter
- |
  draftily
- |
  draftiness
- |
  drafting
- |
  draftsman
- |
  draftswoman
- |
  drafty
- |
  dragger
- |
  draggy
- |
  dragnet
- |
  dragoman
- |
  dragon
- |
  dragonfly
- |
  dragoon
- |
  dragster
- |
  drain
- |
  drainage
- |
  drainboard
- |
  drained
- |
  drainer
- |
  draining
- |
  drainpipe
- |
  Drake
- |
  drake
- |
  Drakensberg
- |
  drama
- |
  Dramamine
- |
  dramatic
- |
  dramatically
- |
  dramatics
- |
  dramatise
- |
  dramatist
- |
  dramatize
- |
  dramaturgic
- |
  dramaturgy
- |
  drank
- |
  drape
- |
  draper
- |
  draperies
- |
  drapery
- |
  drapes
- |
  drastic
- |
  drastically
- |
  draught
- |
  draughts
- |
  draughtsman
- |
  draughty
- |
  Dravidian
- |
  drawback
- |
  drawbridge
- |
  drawee
- |
  drawer
- |
  drawers
- |
  drawing
- |
  drawl
- |
  drawn
- |
  drawstring
- |
  dread
- |
  dreaded
- |
  dreadful
- |
  dreadfully
- |
  dreadfulness
- |
  dreadlocks
- |
  dreadnaught
- |
  dreadnought
- |
  dreads
- |
  dream
- |
  dreamer
- |
  dreamily
- |
  dreaminess
- |
  dreamland
- |
  dreamless
- |
  dreamlike
- |
  dreamt
- |
  dreamworld
- |
  dreamy
- |
  drear
- |
  drearily
- |
  dreariness
- |
  dreary
- |
  dredge
- |
  dredger
- |
  dreggy
- |
  dregs
- |
  dreidel
- |
  dreidl
- |
  Dreiser
- |
  drench
- |
  Dresden
- |
  dress
- |
  dressage
- |
  dressed
- |
  dresser
- |
  dressiness
- |
  dressing
- |
  dressmaker
- |
  dressmaking
- |
  dressy
- |
  Dreyfus
- |
  dribble
- |
  dribbler
- |
  driblet
- |
  dried
- |
  drier
- |
  dries
- |
  driest
- |
  drift
- |
  drifter
- |
  driftwood
- |
  drifty
- |
  drill
- |
  driller
- |
  drilling
- |
  drillmaster
- |
  drily
- |
  drink
- |
  drinkability
- |
  drinkable
- |
  drinker
- |
  drinking
- |
  dripper
- |
  dripping
- |
  drippings
- |
  drivability
- |
  drivable
- |
  drive
- |
  drivel
- |
  driveler
- |
  driveline
- |
  driveller
- |
  driven
- |
  driver
- |
  driveshaft
- |
  drivetrain
- |
  driveway
- |
  driving
- |
  drizzle
- |
  drizzly
- |
  drogue
- |
  droll
- |
  drollery
- |
  drollness
- |
  drolly
- |
  dromedary
- |
  drone
- |
  droning
- |
  drool
- |
  droop
- |
  droopily
- |
  droopiness
- |
  droopingly
- |
  droopy
- |
  dropkick
- |
  droplet
- |
  dropout
- |
  dropper
- |
  dropping
- |
  droppings
- |
  drops
- |
  dropsical
- |
  dropsy
- |
  drosophila
- |
  dross
- |
  drossy
- |
  drought
- |
  drouth
- |
  drove
- |
  drover
- |
  droves
- |
  drown
- |
  drowning
- |
  drowse
- |
  drowsily
- |
  drowsiness
- |
  drowsy
- |
  drubber
- |
  drubbing
- |
  drudge
- |
  drudgery
- |
  druggie
- |
  druggist
- |
  druggy
- |
  drugstore
- |
  Druid
- |
  druid
- |
  Druidic
- |
  druidic
- |
  Druidical
- |
  druidical
- |
  Druidism
- |
  druidism
- |
  drumbeat
- |
  drumlin
- |
  drummer
- |
  drumming
- |
  drumstick
- |
  drunk
- |
  drunkard
- |
  drunken
- |
  drunkenly
- |
  drunkenness
- |
  drupe
- |
  drupelet
- |
  Druse
- |
  Druze
- |
  Dryad
- |
  dryad
- |
  Dryden
- |
  dryer
- |
  dryly
- |
  dryness
- |
  drywall
- |
  Duala
- |
  dualism
- |
  dualist
- |
  dualistic
- |
  duality
- |
  dually
- |
  Duane
- |
  Dubai
- |
  Dubayy
- |
  dubber
- |
  dubbin
- |
  Dubcek
- |
  Dubhe
- |
  dubiety
- |
  dubiosity
- |
  dubious
- |
  dubiously
- |
  dubiousness
- |
  Dublin
- |
  Dubliner
- |
  dubnium
- |
  DuBois
- |
  Dubrovnik
- |
  Dubuque
- |
  ducal
- |
  ducat
- |
  Duchamp
- |
  duchess
- |
  duchy
- |
  duckbill
- |
  duckboard
- |
  duckling
- |
  duckpin
- |
  duckpins
- |
  ducks
- |
  duckweed
- |
  ducky
- |
  ducted
- |
  ductile
- |
  ductility
- |
  ductless
- |
  duded
- |
  dudgeon
- |
  dudish
- |
  Dudley
- |
  dueler
- |
  duelist
- |
  dueller
- |
  duellist
- |
  duende
- |
  duenna
- |
  duffer
- |
  dugout
- |
  Duisburg
- |
  dukedom
- |
  dukes
- |
  dulcet
- |
  dulcify
- |
  dulcimer
- |
  dulcimore
- |
  dullard
- |
  Dulles
- |
  dullish
- |
  dullness
- |
  dully
- |
  dulness
- |
  Duluth
- |
  Dumas
- |
  dumbbell
- |
  dumbfound
- |
  dumbfounded
- |
  dumbly
- |
  dumbness
- |
  dumbwaiter
- |
  dumdum
- |
  dumfound
- |
  Dumfries
- |
  dummy
- |
  dumper
- |
  dumpily
- |
  dumpiness
- |
  dumping
- |
  dumpling
- |
  dumps
- |
  Dumpster
- |
  dumpster
- |
  dumpy
- |
  Dunbar
- |
  Duncan
- |
  dunce
- |
  Dundee
- |
  dunderhead
- |
  Dungannon
- |
  dungaree
- |
  dungarees
- |
  dungeon
- |
  dunghill
- |
  Dunkirk
- |
  dunno
- |
  duodecimal
- |
  duodena
- |
  duodenal
- |
  duodenum
- |
  dupability
- |
  dupable
- |
  duper
- |
  duple
- |
  duplex
- |
  duplicate
- |
  duplication
- |
  duplicator
- |
  duplicitous
- |
  duplicity
- |
  durability
- |
  durable
- |
  durableness
- |
  durably
- |
  durance
- |
  Durango
- |
  Durant
- |
  duration
- |
  Durban
- |
  Durer
- |
  duress
- |
  Durey
- |
  Durga
- |
  Durham
- |
  during
- |
  Durius
- |
  Durkheim
- |
  durrie
- |
  durst
- |
  durum
- |
  Durward
- |
  Dushanbe
- |
  duskiness
- |
  dusky
- |
  Dusseldorf
- |
  dustbin
- |
  duster
- |
  dustiness
- |
  dusting
- |
  dustless
- |
  dustpan
- |
  dusty
- |
  Dutch
- |
  dutch
- |
  Dutchman
- |
  Dutchwoman
- |
  duteous
- |
  duteously
- |
  dutiable
- |
  dutiful
- |
  dutifully
- |
  dutifulness
- |
  Duvalier
- |
  duvet
- |
  Dvorak
- |
  Dwaine
- |
  dwarf
- |
  dwarfed
- |
  dwarfish
- |
  dwarfishness
- |
  dwarfism
- |
  dwarves
- |
  Dwayne
- |
  dweeb
- |
  dwell
- |
  dweller
- |
  dwelling
- |
  dwelt
- |
  Dwight
- |
  dwindle
- |
  dwindling
- |
  dyadic
- |
  dybbuk
- |
  dybbukim
- |
  dyestuff
- |
  Dyfed
- |
  dying
- |
  Dylan
- |
  dynamic
- |
  dynamical
- |
  dynamically
- |
  dynamicist
- |
  dynamics
- |
  dynamism
- |
  dynamist
- |
  dynamite
- |
  dynamo
- |
  dynamometer
- |
  dynamometry
- |
  dynast
- |
  dynastic
- |
  dynastically
- |
  dynasty
- |
  dysenteric
- |
  dysentery
- |
  dysfunction
- |
  dysgenic
- |
  dyslectic
- |
  dyslexia
- |
  dyslexic
- |
  dyspepsia
- |
  dyspeptic
- |
  dysphasia
- |
  dysphasias
- |
  dysphasic
- |
  dysphemism
- |
  dysphoria
- |
  dysphoric
- |
  dysplasia
- |
  dysplastic
- |
  dysprosium
- |
  dystopia
- |
  dystopian
- |
  dystrophic
- |
  dystrophy
- |
  Dzerzhinsk
- |
  Dzerzhinsky
- |
  Eadwig
- |
  eager
- |
  eagerly
- |
  eagerness
- |
  eagle
- |
  eaglet
- |
  Eakins
- |
  Ealing
- |
  earache
- |
  eardrum
- |
  eared
- |
  earflap
- |
  earful
- |
  Earhart
- |
  earldom
- |
  Earle
- |
  earless
- |
  earlier
- |
  earliest
- |
  earliness
- |
  earlobe
- |
  early
- |
  earmark
- |
  earmuff
- |
  earmuffs
- |
  earner
- |
  Earnest
- |
  earnest
- |
  earnestly
- |
  earnestness
- |
  earnings
- |
  earphone
- |
  earphones
- |
  earpiece
- |
  earplug
- |
  earring
- |
  earshot
- |
  earsplitting
- |
  Earth
- |
  earth
- |
  earthbound
- |
  earthed
- |
  earthen
- |
  earthenware
- |
  earthily
- |
  earthiness
- |
  earthliness
- |
  earthling
- |
  earthly
- |
  earthmover
- |
  earthmoving
- |
  earthquake
- |
  earthshaking
- |
  earthward
- |
  earthwards
- |
  earthwork
- |
  earthworm
- |
  earthy
- |
  earwax
- |
  earwig
- |
  easel
- |
  easement
- |
  easily
- |
  easiness
- |
  eastbound
- |
  Easter
- |
  easterly
- |
  Eastern
- |
  eastern
- |
  Easterner
- |
  easterner
- |
  easternmost
- |
  Eastman
- |
  eastward
- |
  eastwardly
- |
  eastwards
- |
  Eastwood
- |
  easygoing
- |
  eatable
- |
  eaten
- |
  eater
- |
  eatery
- |
  eaves
- |
  eavesdrop
- |
  eavesdropper
- |
  EBCDIC
- |
  Ebeneezer
- |
  Eblana
- |
  Ebola
- |
  ebonite
- |
  ebony
- |
  ebullience
- |
  ebulliency
- |
  ebullient
- |
  ebulliently
- |
  ebullition
- |
  eccentric
- |
  eccentricity
- |
  ecclesial
- |
  Ecclesiastes
- |
  ecclesiastic
- |
  ecdyses
- |
  ecdysiasm
- |
  ecdysiast
- |
  ecdysis
- |
  echelon
- |
  echeloning
- |
  echinacea
- |
  echinoderm
- |
  echoer
- |
  echogram
- |
  echoic
- |
  echolalia
- |
  echolocate
- |
  echolocation
- |
  eclair
- |
  eclat
- |
  Eclectic
- |
  eclectic
- |
  eclectically
- |
  eclecticism
- |
  eclipse
- |
  ecliptic
- |
  eclogue
- |
  ecocidal
- |
  ecocide
- |
  ecologic
- |
  ecological
- |
  ecologically
- |
  ecologist
- |
  ecology
- |
  econometric
- |
  econometrics
- |
  econometrist
- |
  economic
- |
  economical
- |
  economically
- |
  economics
- |
  economies
- |
  economism
- |
  economist
- |
  economize
- |
  economizer
- |
  economy
- |
  ecosystem
- |
  ecotourism
- |
  Ecstasy
- |
  ecstasy
- |
  ecstatic
- |
  ecstatically
- |
  ectomorph
- |
  ectomorphic
- |
  ectomorphy
- |
  ectopic
- |
  ectoplasm
- |
  ectoplasmic
- |
  ectotherm
- |
  ectothermal
- |
  ectothermic
- |
  ectothermous
- |
  Ecuador
- |
  Ecuadoran
- |
  Ecuadorean
- |
  Ecuadorian
- |
  ecumenic
- |
  ecumenical
- |
  ecumenically
- |
  ecumenicism
- |
  ecumenism
- |
  ecumenist
- |
  eczema
- |
  eczematous
- |
  edacious
- |
  edacity
- |
  Eddie
- |
  edelweiss
- |
  edema
- |
  edemata
- |
  edematous
- |
  Edenic
- |
  Edgar
- |
  edged
- |
  edger
- |
  edgeways
- |
  edgewise
- |
  edgily
- |
  edginess
- |
  edging
- |
  edibility
- |
  edible
- |
  edibleness
- |
  edict
- |
  edification
- |
  edifice
- |
  edifier
- |
  edify
- |
  Edinburgh
- |
  Edison
- |
  Edith
- |
  edition
- |
  editor
- |
  editorial
- |
  editorialist
- |
  editorialize
- |
  editorially
- |
  editorship
- |
  editress
- |
  Edmond
- |
  Edmonton
- |
  Edmund
- |
  Edomite
- |
  Edson
- |
  educability
- |
  educable
- |
  educate
- |
  educated
- |
  education
- |
  educational
- |
  educative
- |
  educator
- |
  educe
- |
  educible
- |
  eduction
- |
  edutainment
- |
  Edward
- |
  Edwardian
- |
  Edwards
- |
  Edwin
- |
  Edwina
- |
  Edythe
- |
  eerie
- |
  eerily
- |
  eeriness
- |
  efface
- |
  effaceable
- |
  effacement
- |
  effacer
- |
  effect
- |
  effective
- |
  effectively
- |
  effectivity
- |
  effector
- |
  effects
- |
  effectual
- |
  effectuality
- |
  effectually
- |
  effectuate
- |
  effectuation
- |
  effeminacy
- |
  effeminate
- |
  effeminately
- |
  effendi
- |
  efferent
- |
  effervesce
- |
  effervescent
- |
  effete
- |
  effetely
- |
  effeteness
- |
  efficacious
- |
  efficacy
- |
  efficiency
- |
  efficient
- |
  efficiently
- |
  Effie
- |
  effigy
- |
  effleurage
- |
  effloresce
- |
  efflorescent
- |
  effluence
- |
  effluent
- |
  effluvia
- |
  effluvial
- |
  effluvium
- |
  effort
- |
  effortless
- |
  effortlessly
- |
  effrontery
- |
  effulgence
- |
  effulgent
- |
  effulgently
- |
  effuse
- |
  effusion
- |
  effusive
- |
  effusively
- |
  effusiveness
- |
  egads
- |
  egalitarian
- |
  Egbert
- |
  eggbeater
- |
  egghead
- |
  eggnog
- |
  eggplant
- |
  eggshell
- |
  eglantine
- |
  egocentric
- |
  egocentrism
- |
  egoism
- |
  egoist
- |
  egoistic
- |
  egoistical
- |
  egoistically
- |
  egoless
- |
  egomania
- |
  egomaniac
- |
  egomaniacal
- |
  egotism
- |
  egotist
- |
  egotistic
- |
  egotistical
- |
  egotize
- |
  egregious
- |
  egregiously
- |
  egress
- |
  egret
- |
  Egypt
- |
  Egyptian
- |
  Eichmann
- |
  eider
- |
  eiderdown
- |
  eidetic
- |
  eidetically
- |
  eidola
- |
  eidolon
- |
  eidos
- |
  Eiffel
- |
  eight
- |
  eightball
- |
  eighteen
- |
  eighteenth
- |
  eightfold
- |
  eighth
- |
  eightieth
- |
  eighty
- |
  Eileen
- |
  Eindhoven
- |
  Einstein
- |
  einsteinium
- |
  eirenic
- |
  Eisenhower
- |
  Eisenstein
- |
  either
- |
  ejaculate
- |
  ejaculation
- |
  ejaculator
- |
  ejaculatory
- |
  eject
- |
  ejection
- |
  ejector
- |
  elaborate
- |
  elaborately
- |
  elaboration
- |
  elaborative
- |
  elaborator
- |
  Elaine
- |
  Elamite
- |
  eland
- |
  elapid
- |
  elapse
- |
  elasmobranch
- |
  elastic
- |
  elastically
- |
  elasticity
- |
  elasticize
- |
  elate
- |
  elated
- |
  elatedly
- |
  elatedness
- |
  elation
- |
  Elbert
- |
  elbow
- |
  elbowroom
- |
  Elbrus
- |
  Elburz
- |
  elder
- |
  elderberry
- |
  elderly
- |
  eldest
- |
  Eldorado
- |
  eldritch
- |
  Eleanor
- |
  Eleanore
- |
  elect
- |
  electability
- |
  electable
- |
  elected
- |
  election
- |
  electioneer
- |
  elective
- |
  elector
- |
  electoral
- |
  electorally
- |
  electorate
- |
  Electra
- |
  electric
- |
  electrical
- |
  electrically
- |
  electrician
- |
  electricity
- |
  electrified
- |
  electrifier
- |
  electrify
- |
  electrifying
- |
  electrocute
- |
  electrode
- |
  electrolysis
- |
  electrolyte
- |
  electrolytic
- |
  electrolyze
- |
  electron
- |
  electronic
- |
  electronics
- |
  electroplate
- |
  electroscope
- |
  electroshock
- |
  electrotype
- |
  electrotyper
- |
  electrotypic
- |
  eleemosynary
- |
  elegance
- |
  elegant
- |
  elegantly
- |
  elegiac
- |
  elegiacal
- |
  elegiacally
- |
  elegiacs
- |
  elegist
- |
  elegize
- |
  elegy
- |
  element
- |
  elemental
- |
  elementally
- |
  elementarily
- |
  elementary
- |
  elements
- |
  Elena
- |
  elephant
- |
  elephantine
- |
  elevate
- |
  elevation
- |
  elevator
- |
  eleven
- |
  eleventh
- |
  elfin
- |
  elfish
- |
  Elgar
- |
  Elias
- |
  elicit
- |
  elicitation
- |
  elicitor
- |
  elide
- |
  elided
- |
  eligibility
- |
  eligible
- |
  eligibly
- |
  Elijah
- |
  eliminate
- |
  elimination
- |
  eliminative
- |
  eliminator
- |
  eliminatory
- |
  Elinor
- |
  Eliot
- |
  Elisabeth
- |
  Elise
- |
  Elisha
- |
  elision
- |
  elite
- |
  elitism
- |
  elitist
- |
  elixir
- |
  Eliza
- |
  Elizabeth
- |
  Elizabethan
- |
  Ellen
- |
  Ellesmere
- |
  Ellice
- |
  Ellington
- |
  Elliot
- |
  Elliott
- |
  ellipse
- |
  ellipses
- |
  ellipsis
- |
  ellipsoid
- |
  ellipsoidal
- |
  elliptic
- |
  elliptical
- |
  elliptically
- |
  Ellis
- |
  Ellison
- |
  Ellsworth
- |
  Ellwood
- |
  Ellyn
- |
  Elmer
- |
  Elnath
- |
  elocution
- |
  elocutionary
- |
  elocutionist
- |
  elodea
- |
  Eloise
- |
  elongate
- |
  elongated
- |
  elongation
- |
  elope
- |
  elopement
- |
  eloper
- |
  eloquence
- |
  eloquent
- |
  eloquently
- |
  elsewhere
- |
  Elsie
- |
  Elton
- |
  elucidate
- |
  elucidation
- |
  elucidative
- |
  elucidator
- |
  elucidatory
- |
  elude
- |
  eluder
- |
  elusive
- |
  elusively
- |
  elusiveness
- |
  elusory
- |
  elute
- |
  elution
- |
  elver
- |
  elves
- |
  Elvin
- |
  Elvira
- |
  Elwood
- |
  Elysian
- |
  Elysium
- |
  emaciate
- |
  emaciated
- |
  emaciation
- |
  email
- |
  emalangeni
- |
  emanate
- |
  emanation
- |
  emanative
- |
  emanator
- |
  emancipate
- |
  emancipated
- |
  emancipation
- |
  emancipator
- |
  emancipatory
- |
  emasculate
- |
  emasculated
- |
  emasculation
- |
  emasculative
- |
  emasculator
- |
  emasculatory
- |
  embalm
- |
  embalmer
- |
  embalming
- |
  embalmment
- |
  embank
- |
  embankment
- |
  embarcadero
- |
  embargo
- |
  embark
- |
  embarkation
- |
  embarrass
- |
  embarrassed
- |
  embarrassing
- |
  embassy
- |
  embattle
- |
  embattled
- |
  embed
- |
  embedded
- |
  embedment
- |
  embellish
- |
  embellisher
- |
  ember
- |
  embers
- |
  embezzle
- |
  embezzlement
- |
  embezzler
- |
  embitter
- |
  embittered
- |
  embitterment
- |
  emblazon
- |
  emblazoner
- |
  emblazonment
- |
  emblem
- |
  emblematic
- |
  emblematical
- |
  embodiment
- |
  embody
- |
  embolden
- |
  emboli
- |
  embolism
- |
  embolus
- |
  embonpoint
- |
  emboss
- |
  embossed
- |
  embosser
- |
  embossment
- |
  embouchure
- |
  embower
- |
  embrace
- |
  embraceable
- |
  embracement
- |
  embrasure
- |
  embrasured
- |
  embrocate
- |
  embrocation
- |
  embroider
- |
  embroiderer
- |
  embroidery
- |
  embroil
- |
  embroiled
- |
  embroilment
- |
  embrue
- |
  embryo
- |
  embryologic
- |
  embryologist
- |
  embryology
- |
  embryonal
- |
  embryonic
- |
  emcee
- |
  emend
- |
  emendable
- |
  emendation
- |
  emender
- |
  emerald
- |
  emerge
- |
  emergence
- |
  emergency
- |
  emergent
- |
  emerita
- |
  emeritus
- |
  Emerson
- |
  Emersonian
- |
  Emery
- |
  emery
- |
  emetic
- |
  emigrant
- |
  emigrate
- |
  emigration
- |
  emigre
- |
  Emile
- |
  Emilie
- |
  Emily
- |
  eminence
- |
  eminent
- |
  eminently
- |
  emirate
- |
  emissary
- |
  emission
- |
  emitter
- |
  Emmanuel
- |
  Emmet
- |
  emollience
- |
  emollient
- |
  emolument
- |
  emoluments
- |
  Emory
- |
  emote
- |
  emoter
- |
  emoticon
- |
  emotion
- |
  emotional
- |
  emotionalism
- |
  emotionalize
- |
  emotionally
- |
  emotive
- |
  emotively
- |
  emotiveness
- |
  emotivity
- |
  empanada
- |
  empanel
- |
  empathetic
- |
  empathic
- |
  empathically
- |
  empathize
- |
  empathy
- |
  Empedocles
- |
  empennage
- |
  emperor
- |
  emphases
- |
  emphasis
- |
  emphasise
- |
  emphasize
- |
  emphatic
- |
  emphatically
- |
  emphysema
- |
  emphysemic
- |
  empire
- |
  empiric
- |
  empirical
- |
  empirically
- |
  empiricism
- |
  empiricist
- |
  emplacement
- |
  employ
- |
  employable
- |
  employe
- |
  employee
- |
  employer
- |
  employment
- |
  emporia
- |
  emporium
- |
  empower
- |
  empowerment
- |
  empress
- |
  emptily
- |
  emptiness
- |
  empty
- |
  empyreal
- |
  empyrean
- |
  emulate
- |
  emulation
- |
  emulative
- |
  emulator
- |
  emulous
- |
  emulsifier
- |
  emulsify
- |
  emulsion
- |
  emulsive
- |
  enable
- |
  enabler
- |
  enabling
- |
  enact
- |
  enactment
- |
  enactor
- |
  enamel
- |
  enameler
- |
  enameller
- |
  enamelware
- |
  enamor
- |
  enamored
- |
  enamour
- |
  encamp
- |
  encampment
- |
  encapsulate
- |
  encase
- |
  encasement
- |
  enceinte
- |
  encephala
- |
  encephalitic
- |
  encephalitis
- |
  encephalon
- |
  encephalous
- |
  enchain
- |
  enchainment
- |
  enchant
- |
  enchanted
- |
  enchantedly
- |
  enchanter
- |
  enchanting
- |
  enchantingly
- |
  enchantment
- |
  enchantress
- |
  enchilada
- |
  encipher
- |
  encipherment
- |
  encircle
- |
  encirclement
- |
  enclave
- |
  enclitic
- |
  enclitically
- |
  enclose
- |
  enclosed
- |
  enclosure
- |
  encode
- |
  encoder
- |
  encomia
- |
  encomiast
- |
  encomiastic
- |
  encomium
- |
  encompass
- |
  encore
- |
  encounter
- |
  encourage
- |
  encouraged
- |
  encourager
- |
  encouraging
- |
  encroach
- |
  encroacher
- |
  encroachment
- |
  encrust
- |
  encrustation
- |
  encrusted
- |
  encrypt
- |
  encryption
- |
  encumber
- |
  encumbrance
- |
  encyclical
- |
  encyclopedia
- |
  encyclopedic
- |
  encyst
- |
  encystation
- |
  encystment
- |
  endanger
- |
  endangered
- |
  endangerment
- |
  endear
- |
  endearing
- |
  endearingly
- |
  endearment
- |
  endeavor
- |
  endeavour
- |
  Endecott
- |
  endemic
- |
  endemically
- |
  endemicity
- |
  endemism
- |
  Endicott
- |
  ending
- |
  endive
- |
  endless
- |
  endlessly
- |
  endlessness
- |
  endmost
- |
  endnote
- |
  endocrine
- |
  endodontic
- |
  endodontics
- |
  endodontist
- |
  endogamic
- |
  endogamous
- |
  endogamy
- |
  endogenous
- |
  endogenously
- |
  endometria
- |
  endometrial
- |
  endometrium
- |
  endomorph
- |
  endomorphic
- |
  endomorphy
- |
  endoplasm
- |
  endoplasmic
- |
  endorphin
- |
  endorsable
- |
  endorse
- |
  endorsement
- |
  endorser
- |
  endorsor
- |
  endoscope
- |
  endoscopic
- |
  endoscopy
- |
  endotherm
- |
  endothermal
- |
  endothermic
- |
  endow
- |
  endower
- |
  endowment
- |
  endue
- |
  endurable
- |
  endurance
- |
  endure
- |
  enduring
- |
  endways
- |
  endwise
- |
  Endymion
- |
  enema
- |
  enemata
- |
  enemy
- |
  energetic
- |
  energise
- |
  energize
- |
  energizer
- |
  energizing
- |
  energy
- |
  enervate
- |
  enervation
- |
  enervative
- |
  enervator
- |
  Enewetak
- |
  enfeeble
- |
  enfeeblement
- |
  Enfield
- |
  enfilade
- |
  enfold
- |
  enforce
- |
  enforceable
- |
  enforcement
- |
  enforcer
- |
  enfranchise
- |
  engage
- |
  engaged
- |
  engagement
- |
  engager
- |
  engaging
- |
  engagingly
- |
  Engels
- |
  engender
- |
  engine
- |
  engineer
- |
  engineering
- |
  England
- |
  English
- |
  english
- |
  Englishman
- |
  Englishwoman
- |
  Englishwomen
- |
  engorge
- |
  engorged
- |
  engorgement
- |
  engraft
- |
  engram
- |
  engrammatic
- |
  engrave
- |
  engraver
- |
  engraving
- |
  engross
- |
  engrossed
- |
  engrossing
- |
  engrossment
- |
  engulf
- |
  engulfment
- |
  enhance
- |
  enhancement
- |
  enhancer
- |
  enigma
- |
  enigmata
- |
  enigmatic
- |
  enigmatical
- |
  Eniwetok
- |
  enjambement
- |
  enjambment
- |
  enjoin
- |
  enjoinder
- |
  enjoiner
- |
  enjoinment
- |
  enjoy
- |
  enjoyable
- |
  enjoyably
- |
  enjoyer
- |
  enjoyment
- |
  enlarge
- |
  enlargeable
- |
  enlarged
- |
  enlargement
- |
  enlarger
- |
  enlighten
- |
  enlightened
- |
  enlightener
- |
  enlightening
- |
  enlist
- |
  enlisted
- |
  enlistee
- |
  enlistment
- |
  enliven
- |
  enlivenment
- |
  enmesh
- |
  enmeshment
- |
  enmity
- |
  ennead
- |
  Enniskillen
- |
  Ennius
- |
  ennoble
- |
  ennoblement
- |
  ennobling
- |
  ennui
- |
  Enoch
- |
  enologist
- |
  enology
- |
  enormity
- |
  enormous
- |
  enormously
- |
  enormousness
- |
  enough
- |
  enplane
- |
  enquire
- |
  enquirer
- |
  enquiry
- |
  enrage
- |
  enraged
- |
  enrapture
- |
  enrich
- |
  enrichment
- |
  enrol
- |
  enroll
- |
  enrollment
- |
  enrolment
- |
  Enron
- |
  Enschede
- |
  ensconce
- |
  ensemble
- |
  ensheathe
- |
  enshrine
- |
  enshrinement
- |
  enshroud
- |
  ensign
- |
  ensilage
- |
  ensile
- |
  enslave
- |
  enslavement
- |
  enslaver
- |
  ensnare
- |
  ensnarement
- |
  ensnarer
- |
  ensue
- |
  ensuing
- |
  ensure
- |
  ensurer
- |
  entablature
- |
  entail
- |
  entailment
- |
  entangle
- |
  entanglement
- |
  entente
- |
  enter
- |
  enteral
- |
  enteric
- |
  enteritis
- |
  enterprise
- |
  enterprising
- |
  entertain
- |
  entertainer
- |
  entertaining
- |
  enthral
- |
  enthrall
- |
  enthralling
- |
  enthrallment
- |
  enthralment
- |
  enthrone
- |
  enthronement
- |
  enthuse
- |
  enthusiasm
- |
  enthusiast
- |
  enthusiastic
- |
  entice
- |
  enticement
- |
  enticer
- |
  enticing
- |
  enticingly
- |
  entire
- |
  entirely
- |
  entirety
- |
  entitative
- |
  entitle
- |
  entitlement
- |
  entity
- |
  entomb
- |
  entombment
- |
  entomologic
- |
  entomologist
- |
  entomology
- |
  entourage
- |
  entrails
- |
  entrain
- |
  entrance
- |
  entranced
- |
  entrancement
- |
  entrancing
- |
  entrancingly
- |
  entrant
- |
  entrap
- |
  entrapment
- |
  entrapper
- |
  entreat
- |
  entreatingly
- |
  entreatment
- |
  entreaty
- |
  entrechat
- |
  entree
- |
  entrench
- |
  entrenched
- |
  entrenchment
- |
  entrepot
- |
  entrepreneur
- |
  entropic
- |
  entropically
- |
  entropy
- |
  entrust
- |
  entry
- |
  entwine
- |
  enumerable
- |
  enumerate
- |
  enumeration
- |
  enumerative
- |
  enumerator
- |
  enunciate
- |
  enunciation
- |
  enunciative
- |
  enunciator
- |
  enure
- |
  enuresis
- |
  enuretic
- |
  envelop
- |
  envelope
- |
  enveloper
- |
  enveloping
- |
  envelopment
- |
  envenom
- |
  enviability
- |
  enviable
- |
  enviably
- |
  envier
- |
  envious
- |
  enviously
- |
  enviousness
- |
  environment
- |
  environs
- |
  envisage
- |
  envision
- |
  envoi
- |
  envoy
- |
  envyingly
- |
  enzymatic
- |
  enzyme
- |
  enzymic
- |
  enzymically
- |
  Eocene
- |
  eolian
- |
  eonian
- |
  eosin
- |
  epaulet
- |
  epaulette
- |
  ephebe
- |
  ephebic
- |
  ephedrine
- |
  ephemera
- |
  ephemeral
- |
  ephemerality
- |
  ephemerally
- |
  ephemeron
- |
  Ephesian
- |
  Ephesians
- |
  Ephesus
- |
  Ephraim
- |
  Ephraimite
- |
  epical
- |
  epically
- |
  epicene
- |
  epicenter
- |
  epicentral
- |
  Epictetus
- |
  epicure
- |
  Epicurean
- |
  epicurean
- |
  Epicureanism
- |
  epicurism
- |
  Epicurus
- |
  epidemic
- |
  epidemically
- |
  epidemiology
- |
  epidermal
- |
  epidermic
- |
  epidermis
- |
  epidermoid
- |
  epidural
- |
  epiglottal
- |
  epiglottis
- |
  epigram
- |
  epigrammatic
- |
  epigraph
- |
  epigrapher
- |
  epigraphic
- |
  epigraphy
- |
  epilepsy
- |
  epileptic
- |
  epilog
- |
  epilogue
- |
  epinephrin
- |
  epinephrine
- |
  epiphanic
- |
  Epiphany
- |
  epiphany
- |
  epiphytal
- |
  epiphyte
- |
  epiphytic
- |
  episcopacy
- |
  Episcopal
- |
  episcopal
- |
  Episcopalian
- |
  episcopalian
- |
  episcopate
- |
  episiotomy
- |
  episode
- |
  episodic
- |
  episodically
- |
  epistemic
- |
  epistemology
- |
  Epistle
- |
  epistle
- |
  epistolary
- |
  epitaph
- |
  epithalamia
- |
  epithalamion
- |
  epithalamium
- |
  epithelia
- |
  epithelial
- |
  epithelium
- |
  epithet
- |
  epithetic
- |
  epithetical
- |
  epitome
- |
  epitomise
- |
  epitomist
- |
  epitomize
- |
  epoch
- |
  epochal
- |
  epode
- |
  eponym
- |
  eponymous
- |
  epoxy
- |
  epsilon
- |
  equability
- |
  equable
- |
  equably
- |
  equal
- |
  equalise
- |
  equaliser
- |
  equality
- |
  equalization
- |
  equalize
- |
  equalizer
- |
  equally
- |
  equanimity
- |
  equanimous
- |
  equatable
- |
  equate
- |
  equation
- |
  equator
- |
  equatorial
- |
  equerry
- |
  equestrian
- |
  equestrienne
- |
  equiangular
- |
  equidistance
- |
  equidistant
- |
  equilateral
- |
  equilibrate
- |
  equilibria
- |
  equilibrial
- |
  equilibrium
- |
  equine
- |
  equinoctial
- |
  equinox
- |
  equip
- |
  equipage
- |
  equipment
- |
  equipoise
- |
  equipped
- |
  equitability
- |
  equitable
- |
  equitably
- |
  equitation
- |
  equities
- |
  Equity
- |
  equity
- |
  equivalence
- |
  equivalency
- |
  equivalent
- |
  equivalently
- |
  equivocal
- |
  equivocality
- |
  equivocally
- |
  equivocate
- |
  equivocation
- |
  equivocator
- |
  equivocatory
- |
  Equuleus
- |
  eradicable
- |
  eradicant
- |
  eradicate
- |
  eradication
- |
  eradicator
- |
  erasable
- |
  erase
- |
  eraser
- |
  Erasmus
- |
  erasure
- |
  Erbil
- |
  erbium
- |
  Erebus
- |
  erect
- |
  erectile
- |
  erection
- |
  erectly
- |
  erectness
- |
  erector
- |
  erelong
- |
  eremite
- |
  eremitic
- |
  eremitical
- |
  Erevan
- |
  Erfurt
- |
  ergative
- |
  ergativity
- |
  ergonometric
- |
  ergonomic
- |
  ergonomics
- |
  ergonomist
- |
  ergosterol
- |
  ergot
- |
  Erica
- |
  Erich
- |
  Ericson
- |
  Ericsson
- |
  Eridanus
- |
  Erika
- |
  Eriksson
- |
  Eritrea
- |
  Eritrean
- |
  ermine
- |
  Ernest
- |
  Ernestine
- |
  Ernie
- |
  Ernst
- |
  erode
- |
  eroded
- |
  erodible
- |
  erogenic
- |
  erogenous
- |
  erosion
- |
  erosional
- |
  erosionally
- |
  erosive
- |
  erosiveness
- |
  erotic
- |
  erotica
- |
  erotically
- |
  eroticism
- |
  eroticist
- |
  errancy
- |
  errand
- |
  errant
- |
  errantly
- |
  errantry
- |
  errata
- |
  erratic
- |
  erratically
- |
  erraticism
- |
  erratum
- |
  Errol
- |
  erroneous
- |
  erroneously
- |
  error
- |
  errorless
- |
  ersatz
- |
  erstwhile
- |
  eruct
- |
  eructation
- |
  erudite
- |
  eruditely
- |
  erudition
- |
  erupt
- |
  eruption
- |
  eruptive
- |
  Erwin
- |
  erysipelas
- |
  erythema
- |
  erythrocyte
- |
  erythrocytic
- |
  erythromycin
- |
  Erzgebirge
- |
  escalate
- |
  escalation
- |
  escalator
- |
  escallop
- |
  escalop
- |
  escapade
- |
  escape
- |
  escaped
- |
  escapee
- |
  escapement
- |
  escaper
- |
  escapism
- |
  escapist
- |
  escarole
- |
  escarpment
- |
  eschatology
- |
  escheat
- |
  escheated
- |
  Escher
- |
  eschew
- |
  eschewal
- |
  Escondido
- |
  escort
- |
  escritoire
- |
  escrow
- |
  escudo
- |
  esculent
- |
  escutcheon
- |
  escutcheoned
- |
  Esdras
- |
  Esfahan
- |
  Eskimo
- |
  Eskimoan
- |
  Eskisehir
- |
  esophageal
- |
  esophagi
- |
  esophagus
- |
  esoteric
- |
  esoterica
- |
  esoterically
- |
  esotericism
- |
  esotericist
- |
  espadrille
- |
  espalier
- |
  especial
- |
  especially
- |
  Esperantist
- |
  Esperanto
- |
  espionage
- |
  esplanade
- |
  Espoo
- |
  espousal
- |
  espouse
- |
  espouser
- |
  espresso
- |
  esprit
- |
  Esquire
- |
  esquire
- |
  essay
- |
  essayer
- |
  essayist
- |
  Essen
- |
  essence
- |
  Essene
- |
  essential
- |
  essentialism
- |
  essentialist
- |
  essentiality
- |
  essentialize
- |
  essentially
- |
  Essex
- |
  establish
- |
  established
- |
  establisher
- |
  estate
- |
  esteem
- |
  esteemed
- |
  Estella
- |
  Estelle
- |
  ester
- |
  Esther
- |
  esthesia
- |
  esthete
- |
  esthetic
- |
  esthetically
- |
  esthetician
- |
  estheticism
- |
  esthetics
- |
  estimable
- |
  estimably
- |
  estimate
- |
  estimated
- |
  estimation
- |
  estimator
- |
  estival
- |
  estivate
- |
  estivation
- |
  Estonia
- |
  Estonian
- |
  estop
- |
  estoppel
- |
  estrange
- |
  estranged
- |
  estrangement
- |
  estrogen
- |
  estrogenic
- |
  estrous
- |
  estrum
- |
  estrus
- |
  estuarial
- |
  estuarine
- |
  estuary
- |
  etagere
- |
  etcher
- |
  etching
- |
  eternal
- |
  eternally
- |
  eternalness
- |
  eternity
- |
  Ethan
- |
  ethane
- |
  ethanol
- |
  Ethel
- |
  Ethelbert
- |
  Ethelred
- |
  ether
- |
  ethereal
- |
  ethereality
- |
  etherealize
- |
  ethereally
- |
  etherealness
- |
  Ethernet
- |
  ethic
- |
  ethical
- |
  ethically
- |
  ethicist
- |
  ethics
- |
  Ethiopia
- |
  Ethiopian
- |
  ethnic
- |
  ethnically
- |
  ethnicity
- |
  ethnocentric
- |
  ethnographer
- |
  ethnographic
- |
  ethnography
- |
  ethnologic
- |
  ethnological
- |
  ethnologist
- |
  ethnology
- |
  ethological
- |
  ethologist
- |
  ethology
- |
  ethos
- |
  ethyl
- |
  ethylene
- |
  ethyne
- |
  etiologic
- |
  etiological
- |
  etiologist
- |
  etiology
- |
  etiquette
- |
  Etobicoke
- |
  Etruria
- |
  Etrurian
- |
  Etruscan
- |
  etude
- |
  etymological
- |
  etymologist
- |
  etymology
- |
  eucalypti
- |
  eucalyptus
- |
  eucaryote
- |
  Eucharist
- |
  Eucharistic
- |
  eucharistic
- |
  euchre
- |
  Euclid
- |
  Euclidean
- |
  euclidean
- |
  Euclidian
- |
  euclidian
- |
  Eugene
- |
  Eugenia
- |
  eugenic
- |
  eugenically
- |
  eugenicist
- |
  eugenics
- |
  Eugenie
- |
  eugenist
- |
  eukaryote
- |
  eukaryotic
- |
  eulogist
- |
  eulogistic
- |
  eulogize
- |
  eulogizer
- |
  eulogy
- |
  Eunice
- |
  eunuch
- |
  euphemism
- |
  euphemist
- |
  euphemistic
- |
  euphemize
- |
  euphonic
- |
  euphonious
- |
  euphoniously
- |
  euphonize
- |
  euphony
- |
  euphoria
- |
  euphoriant
- |
  euphoric
- |
  Euphrates
- |
  euphuism
- |
  euphuist
- |
  euphuistic
- |
  Eurasia
- |
  Eurasian
- |
  eureka
- |
  Euripidean
- |
  Euripides
- |
  Eurobond
- |
  Eurocentric
- |
  Eurocentrism
- |
  Eurocentrist
- |
  Eurocurrency
- |
  Eurodollar
- |
  Europa
- |
  Europe
- |
  European
- |
  europium
- |
  Eurydice
- |
  eurythmics
- |
  eustacy
- |
  eustasy
- |
  eustatic
- |
  euthanasia
- |
  euthanize
- |
  euthenics
- |
  euthenist
- |
  eutrophic
- |
  eutrophicate
- |
  evacuate
- |
  evacuation
- |
  evacuee
- |
  evade
- |
  evader
- |
  evaluate
- |
  evaluation
- |
  evaluator
- |
  evanesce
- |
  evanescence
- |
  evanescent
- |
  evanescently
- |
  evangelic
- |
  Evangelical
- |
  evangelical
- |
  Evangeline
- |
  evangelism
- |
  Evangelist
- |
  evangelist
- |
  evangelistic
- |
  evangelize
- |
  evangelizer
- |
  Evans
- |
  Evanston
- |
  Evansville
- |
  evaporable
- |
  evaporate
- |
  evaporation
- |
  evaporative
- |
  evaporator
- |
  evaporite
- |
  evasion
- |
  evasive
- |
  evasively
- |
  evasiveness
- |
  Evelyn
- |
  evenhanded
- |
  evenhandedly
- |
  evening
- |
  evenly
- |
  evenness
- |
  evensong
- |
  event
- |
  eventful
- |
  eventfully
- |
  eventfulness
- |
  eventide
- |
  eventual
- |
  eventuality
- |
  eventually
- |
  eventuate
- |
  eventuation
- |
  Everest
- |
  Everett
- |
  everglade
- |
  Everglades
- |
  evergreen
- |
  everlasting
- |
  evermore
- |
  every
- |
  everybody
- |
  everyday
- |
  everyone
- |
  everyplace
- |
  everything
- |
  everywhere
- |
  evict
- |
  eviction
- |
  evictor
- |
  evidence
- |
  evident
- |
  evidential
- |
  evidently
- |
  evildoer
- |
  evildoing
- |
  evilly
- |
  evilness
- |
  evince
- |
  evincible
- |
  eviscerate
- |
  evisceration
- |
  evitable
- |
  evocable
- |
  evocation
- |
  evocative
- |
  evocatively
- |
  evoke
- |
  evoker
- |
  evolution
- |
  evolutionary
- |
  evolutionism
- |
  evolutionist
- |
  evolvable
- |
  evolve
- |
  evolvement
- |
  evulsion
- |
  exacerbate
- |
  exacerbation
- |
  exact
- |
  exactable
- |
  exacting
- |
  exactingly
- |
  exaction
- |
  exactitude
- |
  exactly
- |
  exactness
- |
  exactor
- |
  exaggerate
- |
  exaggerated
- |
  exaggeration
- |
  exaggerative
- |
  exaggerator
- |
  exaggeratory
- |
  exalt
- |
  exaltation
- |
  exalted
- |
  examen
- |
  examination
- |
  examine
- |
  examinee
- |
  examiner
- |
  example
- |
  exasperate
- |
  exasperated
- |
  exasperating
- |
  exasperation
- |
  Excalibur
- |
  excavate
- |
  excavation
- |
  excavator
- |
  exceed
- |
  exceeding
- |
  exceedingly
- |
  excel
- |
  Excellence
- |
  excellence
- |
  Excellency
- |
  excellency
- |
  excellent
- |
  excellently
- |
  excelsior
- |
  except
- |
  excepted
- |
  excepting
- |
  exception
- |
  exceptional
- |
  excerpt
- |
  excess
- |
  excesses
- |
  excessive
- |
  excessively
- |
  exchange
- |
  exchangeable
- |
  Exchequer
- |
  exchequer
- |
  excipient
- |
  excise
- |
  excision
- |
  excitability
- |
  excitable
- |
  excitably
- |
  excitant
- |
  excitation
- |
  excite
- |
  excited
- |
  excitedly
- |
  excitement
- |
  exciter
- |
  exciting
- |
  excitingly
- |
  exclaim
- |
  exclamation
- |
  exclamatory
- |
  exclude
- |
  excluding
- |
  exclusion
- |
  exclusive
- |
  exclusively
- |
  exclusivity
- |
  excogitate
- |
  excoriate
- |
  excoriation
- |
  excrement
- |
  excremental
- |
  excrescence
- |
  excrescent
- |
  excreta
- |
  excrete
- |
  excretion
- |
  excretive
- |
  excretory
- |
  excruciating
- |
  exculpate
- |
  exculpation
- |
  exculpatory
- |
  excursion
- |
  excursionist
- |
  excursive
- |
  excursively
- |
  excursus
- |
  excusable
- |
  excuse
- |
  excuser
- |
  execrable
- |
  execrably
- |
  execrate
- |
  execration
- |
  execrative
- |
  execrator
- |
  execratory
- |
  executable
- |
  execute
- |
  executer
- |
  execution
- |
  executioner
- |
  executive
- |
  executor
- |
  executorial
- |
  executorship
- |
  executory
- |
  executrices
- |
  executrix
- |
  exegeses
- |
  exegesis
- |
  exegete
- |
  exegetic
- |
  exegetical
- |
  exempla
- |
  exemplar
- |
  exemplarily
- |
  exemplarity
- |
  exemplary
- |
  exemplifier
- |
  exemplify
- |
  exemplum
- |
  exempt
- |
  exemptible
- |
  exemption
- |
  exequy
- |
  exercise
- |
  exerciser
- |
  exercises
- |
  exert
- |
  exertion
- |
  Exeter
- |
  exfoliant
- |
  exfoliate
- |
  exfoliation
- |
  exfoliative
- |
  exfoliator
- |
  exhalation
- |
  exhale
- |
  exhaust
- |
  exhausted
- |
  exhaustible
- |
  exhausting
- |
  exhaustion
- |
  exhaustive
- |
  exhaustively
- |
  exhibit
- |
  exhibition
- |
  exhibitor
- |
  exhilarate
- |
  exhilarated
- |
  exhilarating
- |
  exhilaration
- |
  exhilirative
- |
  exhort
- |
  exhortation
- |
  exhortative
- |
  exhortatory
- |
  exhorter
- |
  exhumation
- |
  exhume
- |
  exigence
- |
  exigencies
- |
  exigency
- |
  exigent
- |
  exiguity
- |
  exiguous
- |
  exiguously
- |
  exiguousness
- |
  exile
- |
  exiled
- |
  exist
- |
  existence
- |
  existent
- |
  existential
- |
  existing
- |
  exobiologist
- |
  exobiology
- |
  exocrine
- |
  Exodus
- |
  exodus
- |
  exogamous
- |
  exogamy
- |
  exogenous
- |
  exogenously
- |
  exonerate
- |
  exoneration
- |
  exonerative
- |
  exonerator
- |
  exorbitance
- |
  exorbitant
- |
  exorbitantly
- |
  exorcise
- |
  exorcism
- |
  exorcist
- |
  exorcize
- |
  exoskeletal
- |
  exoskeleton
- |
  exosphere
- |
  exospheric
- |
  exoteric
- |
  exothermal
- |
  exothermic
- |
  exotic
- |
  exotically
- |
  exoticism
- |
  expand
- |
  expandable
- |
  expander
- |
  expanse
- |
  expansible
- |
  expansion
- |
  expansionary
- |
  expansionism
- |
  expansionist
- |
  expansive
- |
  expansively
- |
  expatiate
- |
  expatiation
- |
  expatriate
- |
  expatriation
- |
  expect
- |
  expectancy
- |
  expectant
- |
  expectantly
- |
  expectation
- |
  expectations
- |
  expectorant
- |
  expectorate
- |
  expedience
- |
  expediency
- |
  expedient
- |
  expediently
- |
  expedite
- |
  expediter
- |
  expedition
- |
  expeditious
- |
  expeditor
- |
  expel
- |
  expellable
- |
  expeller
- |
  expend
- |
  expendable
- |
  expender
- |
  expenditure
- |
  expense
- |
  expenses
- |
  expensive
- |
  expensively
- |
  experience
- |
  experienced
- |
  experiential
- |
  experiment
- |
  experimental
- |
  experimenter
- |
  expert
- |
  expertise
- |
  expertly
- |
  expertness
- |
  expiable
- |
  expiate
- |
  expiation
- |
  expiator
- |
  expiatory
- |
  expiration
- |
  expire
- |
  expiry
- |
  explain
- |
  explainable
- |
  explainer
- |
  explanation
- |
  explanatory
- |
  expletive
- |
  explicable
- |
  explicably
- |
  explicate
- |
  explication
- |
  explicative
- |
  explicator
- |
  explicatory
- |
  explicit
- |
  explicitly
- |
  explicitness
- |
  explodable
- |
  explode
- |
  exploded
- |
  exploder
- |
  exploit
- |
  exploitable
- |
  exploitation
- |
  exploitative
- |
  exploiter
- |
  exploitive
- |
  exploration
- |
  exploratory
- |
  explore
- |
  explorer
- |
  explosion
- |
  explosive
- |
  explosively
- |
  exponent
- |
  exponential
- |
  export
- |
  exportable
- |
  exportation
- |
  exporter
- |
  expose
- |
  exposed
- |
  exposer
- |
  exposition
- |
  expositional
- |
  expositor
- |
  expository
- |
  expostulate
- |
  expostulator
- |
  exposure
- |
  expound
- |
  expounder
- |
  express
- |
  expressible
- |
  expression
- |
  expressive
- |
  expressively
- |
  expressly
- |
  expressway
- |
  expropriate
- |
  expropriator
- |
  expulsion
- |
  expunction
- |
  expunge
- |
  expungement
- |
  expunger
- |
  expurgate
- |
  expurgated
- |
  expurgation
- |
  expurgator
- |
  expurgatory
- |
  exquisite
- |
  exquisitely
- |
  extant
- |
  extemporary
- |
  extempore
- |
  extemporize
- |
  extend
- |
  extendable
- |
  extended
- |
  extender
- |
  extendible
- |
  extensible
- |
  extension
- |
  extensive
- |
  extensively
- |
  extensor
- |
  extent
- |
  extenuate
- |
  extenuated
- |
  extenuating
- |
  extenuation
- |
  extenuator
- |
  extenuatory
- |
  exterior
- |
  exteriorly
- |
  exterminate
- |
  exterminator
- |
  external
- |
  externalize
- |
  externally
- |
  externals
- |
  extinct
- |
  extinction
- |
  extinguish
- |
  extinguisher
- |
  extirpate
- |
  extirpation
- |
  extirpative
- |
  extirpator
- |
  extol
- |
  extoll
- |
  extoller
- |
  extolment
- |
  extort
- |
  extorter
- |
  extortion
- |
  extortionate
- |
  extortioner
- |
  extortionist
- |
  extortive
- |
  extra
- |
  extract
- |
  extractable
- |
  extractible
- |
  extraction
- |
  extractor
- |
  extraditable
- |
  extradite
- |
  extradition
- |
  extrados
- |
  extralegal
- |
  extralegally
- |
  extramarital
- |
  extramural
- |
  extraneous
- |
  extraneously
- |
  extrapolate
- |
  extrapolated
- |
  extrapolator
- |
  extrasensory
- |
  extravagance
- |
  extravagant
- |
  extravaganza
- |
  extraversion
- |
  extravert
- |
  extraverted
- |
  extreme
- |
  extremely
- |
  extremeness
- |
  extremism
- |
  extremist
- |
  extremities
- |
  extremity
- |
  extricable
- |
  extricate
- |
  extrication
- |
  extrinsic
- |
  extroversion
- |
  extrovert
- |
  extroverted
- |
  extrudable
- |
  extrude
- |
  extruder
- |
  extrusile
- |
  extrusion
- |
  extrusive
- |
  exuberance
- |
  exuberant
- |
  exuberantly
- |
  exudate
- |
  exudation
- |
  exudative
- |
  exude
- |
  exult
- |
  exultant
- |
  exultantly
- |
  exultation
- |
  exultingly
- |
  exurb
- |
  exurban
- |
  exurbanite
- |
  exurbia
- |
  eyeball
- |
  eyebrow
- |
  eyedropper
- |
  eyeful
- |
  eyeglass
- |
  eyeglasses
- |
  eyelash
- |
  eyeless
- |
  eyelet
- |
  eyelid
- |
  eyeliner
- |
  eyeopener
- |
  eyeopening
- |
  eyepiece
- |
  eyeshadow
- |
  eyesight
- |
  eyesore
- |
  eyestrain
- |
  eyeteeth
- |
  eyetooth
- |
  eyewash
- |
  eyewitness
- |
  eyrie
- |
  eyrir
- |
  Eysenck
- |
  Ezechiel
- |
  Ezekiel
- |
  Faberge
- |
  Fabian
- |
  Fabianism
- |
  fable
- |
  fabled
- |
  fabliau
- |
  fabliaux
- |
  fabric
- |
  fabricate
- |
  fabrication
- |
  fabricator
- |
  fabulist
- |
  fabulous
- |
  fabulously
- |
  fabulousness
- |
  facade
- |
  faced
- |
  facedown
- |
  faceless
- |
  facelift
- |
  facet
- |
  faceted
- |
  facetiae
- |
  facetious
- |
  facetiously
- |
  facia
- |
  faciae
- |
  facial
- |
  facially
- |
  facile
- |
  facilely
- |
  facileness
- |
  facilitate
- |
  facilitation
- |
  facilitative
- |
  facilitator
- |
  facilitatory
- |
  facilities
- |
  facility
- |
  facing
- |
  facsimile
- |
  faction
- |
  factional
- |
  factionalism
- |
  factious
- |
  factiously
- |
  factiousness
- |
  factitious
- |
  factitiously
- |
  factoid
- |
  factor
- |
  factorial
- |
  factory
- |
  factotum
- |
  factual
- |
  factuality
- |
  factually
- |
  faculty
- |
  faddish
- |
  faddist
- |
  faded
- |
  fadeout
- |
  faecal
- |
  faeces
- |
  faerie
- |
  Faeroe
- |
  Faeroese
- |
  faery
- |
  faggot
- |
  faggoting
- |
  Fagin
- |
  fagot
- |
  fagoting
- |
  Fahrenheit
- |
  faience
- |
  failing
- |
  faille
- |
  failure
- |
  faineant
- |
  faint
- |
  fainthearted
- |
  faintly
- |
  faintness
- |
  Fairbanks
- |
  Fairfield
- |
  fairground
- |
  fairgrounds
- |
  fairing
- |
  fairly
- |
  fairness
- |
  fairway
- |
  fairy
- |
  fairyland
- |
  fairytale
- |
  Faisal
- |
  Faisalabad
- |
  Faith
- |
  faith
- |
  faithful
- |
  faithfully
- |
  faithfulness
- |
  faithless
- |
  faithlessly
- |
  fajita
- |
  fajitas
- |
  faker
- |
  fakery
- |
  fakir
- |
  falafel
- |
  falcon
- |
  falconer
- |
  falconry
- |
  Falkland
- |
  Falla
- |
  fallacious
- |
  fallaciously
- |
  fallacy
- |
  fallback
- |
  fallen
- |
  fallibility
- |
  fallible
- |
  fallibleness
- |
  fallibly
- |
  falloff
- |
  fallout
- |
  fallow
- |
  fallowness
- |
  falls
- |
  false
- |
  falsehood
- |
  falsely
- |
  falseness
- |
  falsetto
- |
  falsie
- |
  falsifier
- |
  falsify
- |
  falsity
- |
  Falstaff
- |
  falter
- |
  falterer
- |
  faltering
- |
  falteringly
- |
  Falwell
- |
  famed
- |
  familial
- |
  familiar
- |
  familiarity
- |
  familiarize
- |
  familiarly
- |
  family
- |
  famine
- |
  famish
- |
  famished
- |
  famous
- |
  famously
- |
  fanatic
- |
  fanatical
- |
  fanatically
- |
  fanaticism
- |
  fancier
- |
  fanciful
- |
  fancifully
- |
  fancifulness
- |
  fancily
- |
  fanciness
- |
  fancy
- |
  fancywork
- |
  fandango
- |
  fandom
- |
  fanfare
- |
  fanfaronade
- |
  fanged
- |
  fanjet
- |
  fanlight
- |
  Fannie
- |
  Fanny
- |
  fanny
- |
  fantail
- |
  fantailed
- |
  fantasia
- |
  fantasise
- |
  fantasize
- |
  fantasizer
- |
  fantastic
- |
  fantastical
- |
  fantasy
- |
  fanzine
- |
  faquir
- |
  farad
- |
  Faraday
- |
  faraway
- |
  farce
- |
  farceur
- |
  farcical
- |
  farcicality
- |
  farcically
- |
  farer
- |
  farewell
- |
  farfetched
- |
  Fargo
- |
  Faridabad
- |
  farina
- |
  farinaceous
- |
  farmable
- |
  Farmer
- |
  farmer
- |
  farmhand
- |
  farmhouse
- |
  farming
- |
  farmland
- |
  farmstead
- |
  farmyard
- |
  Faroe
- |
  farouche
- |
  Farouk
- |
  farraginous
- |
  farrago
- |
  Farragut
- |
  Farrell
- |
  farrier
- |
  farriery
- |
  farrow
- |
  farseeing
- |
  farsighted
- |
  farther
- |
  farthermost
- |
  farthest
- |
  farthing
- |
  farthingale
- |
  fasces
- |
  fascia
- |
  fasciae
- |
  fascicle
- |
  fascicled
- |
  fascicule
- |
  fasciculus
- |
  fascinate
- |
  fascinated
- |
  fascinating
- |
  fascination
- |
  fascinator
- |
  Fascism
- |
  fascism
- |
  Fascist
- |
  fascist
- |
  Fascistic
- |
  fascistic
- |
  fashion
- |
  fashionable
- |
  fashionably
- |
  fashioner
- |
  Fassbinder
- |
  fastback
- |
  fastball
- |
  fasten
- |
  fastener
- |
  fastening
- |
  fastidious
- |
  fastidiously
- |
  fastigiate
- |
  fasting
- |
  fastness
- |
  fatal
- |
  fatalism
- |
  fatalist
- |
  fatalistic
- |
  fatality
- |
  fatally
- |
  fatback
- |
  fated
- |
  fateful
- |
  fatefully
- |
  fatefulness
- |
  Fates
- |
  fathead
- |
  fatheaded
- |
  Father
- |
  father
- |
  fatherhood
- |
  fatherland
- |
  fatherless
- |
  fatherliness
- |
  fatherly
- |
  fathom
- |
  fathomable
- |
  fathomless
- |
  fatigable
- |
  fatigue
- |
  fatigues
- |
  Fatima
- |
  fatless
- |
  fatly
- |
  fatness
- |
  fatten
- |
  fattener
- |
  fattening
- |
  fattiness
- |
  fattish
- |
  fatty
- |
  fatuity
- |
  fatuous
- |
  fatuously
- |
  fatuousness
- |
  fatwa
- |
  faubourg
- |
  fauces
- |
  faucet
- |
  Faulkner
- |
  Faulknerian
- |
  fault
- |
  faultfinder
- |
  faultfinding
- |
  faultily
- |
  faultiness
- |
  faultless
- |
  faultlessly
- |
  faulty
- |
  fauna
- |
  faunae
- |
  faunal
- |
  faunally
- |
  faunistic
- |
  Faure
- |
  Faust
- |
  Faustian
- |
  Faustus
- |
  Fauve
- |
  fauve
- |
  Fauvism
- |
  fauvism
- |
  Fauvist
- |
  fauvist
- |
  favor
- |
  favorable
- |
  favorably
- |
  favored
- |
  favorer
- |
  favorite
- |
  favoritism
- |
  favors
- |
  favour
- |
  favourable
- |
  favourably
- |
  favoured
- |
  favourite
- |
  Fawkes
- |
  fawner
- |
  fawningly
- |
  Fayetteville
- |
  fealty
- |
  fearer
- |
  fearful
- |
  fearfully
- |
  fearfulness
- |
  fearless
- |
  fearlessly
- |
  fearlessness
- |
  fearsome
- |
  fearsomely
- |
  fearsomeness
- |
  feasibility
- |
  feasible
- |
  feasibleness
- |
  feasibly
- |
  feast
- |
  feaster
- |
  feasting
- |
  feather
- |
  featherbed
- |
  featherbrain
- |
  feathered
- |
  featheredge
- |
  feathering
- |
  featherless
- |
  feathers
- |
  feathery
- |
  feature
- |
  featureless
- |
  features
- |
  feaze
- |
  febrifugal
- |
  febrifuge
- |
  febrile
- |
  febrility
- |
  February
- |
  fecal
- |
  feces
- |
  feckless
- |
  fecklessly
- |
  fecklessness
- |
  feculence
- |
  feculent
- |
  fecund
- |
  fecundate
- |
  fecundation
- |
  fecundity
- |
  fedayeen
- |
  Federal
- |
  federal
- |
  Federalism
- |
  federalism
- |
  Federalist
- |
  federalist
- |
  federalize
- |
  federally
- |
  federate
- |
  federated
- |
  federation
- |
  federative
- |
  federatively
- |
  fedora
- |
  feeble
- |
  feebleminded
- |
  feebleness
- |
  feebly
- |
  feedback
- |
  feedbag
- |
  feeder
- |
  feeding
- |
  feedlot
- |
  feedstock
- |
  feedstuff
- |
  feeler
- |
  feeling
- |
  feelingly
- |
  feelings
- |
  feign
- |
  feigner
- |
  feint
- |
  feistily
- |
  feistiness
- |
  feisty
- |
  felafel
- |
  feldspar
- |
  Felice
- |
  Felicia
- |
  felicitate
- |
  felicitation
- |
  felicitator
- |
  felicitous
- |
  felicitously
- |
  felicity
- |
  feline
- |
  felinity
- |
  Felix
- |
  fella
- |
  fellable
- |
  fellah
- |
  fellaheen
- |
  fellahin
- |
  fellatio
- |
  fellation
- |
  fellator
- |
  feller
- |
  Fellini
- |
  fellow
- |
  fellowman
- |
  fellowship
- |
  felon
- |
  felonious
- |
  felony
- |
  female
- |
  femaleness
- |
  feminine
- |
  femininely
- |
  feminineness
- |
  femininity
- |
  feminism
- |
  feminist
- |
  feminization
- |
  feminize
- |
  femora
- |
  femoral
- |
  femur
- |
  fence
- |
  fencer
- |
  fencing
- |
  fender
- |
  fenestration
- |
  Fenian
- |
  Fenianism
- |
  fennel
- |
  fenny
- |
  feral
- |
  Ferber
- |
  Ferdinand
- |
  Fermanagh
- |
  ferment
- |
  fermentable
- |
  fermentation
- |
  fermentative
- |
  fermented
- |
  Fermi
- |
  fermion
- |
  fermium
- |
  Fernando
- |
  Ferne
- |
  fernery
- |
  ferny
- |
  ferocious
- |
  ferociously
- |
  ferocity
- |
  Ferrara
- |
  Ferraro
- |
  ferret
- |
  ferric
- |
  ferromagnet
- |
  ferrotype
- |
  ferrous
- |
  ferrule
- |
  ferry
- |
  ferryboat
- |
  fertile
- |
  fertilely
- |
  fertileness
- |
  fertilise
- |
  fertiliser
- |
  fertility
- |
  fertilizable
- |
  fertilize
- |
  fertilizer
- |
  ferule
- |
  fervency
- |
  fervent
- |
  fervently
- |
  fervid
- |
  fervidly
- |
  fervidness
- |
  fervor
- |
  fervour
- |
  fescue
- |
  festal
- |
  festally
- |
  fester
- |
  festering
- |
  festival
- |
  festive
- |
  festively
- |
  festiveness
- |
  festivities
- |
  festivity
- |
  festoon
- |
  fetal
- |
  fetch
- |
  fetcher
- |
  fetching
- |
  fetchingly
- |
  fetich
- |
  feticide
- |
  fetid
- |
  fetidly
- |
  fetidness
- |
  fetish
- |
  fetishism
- |
  fetishist
- |
  fetishistic
- |
  fetlock
- |
  fetoscope
- |
  fetter
- |
  fetters
- |
  fettle
- |
  fettuccine
- |
  fetus
- |
  feudal
- |
  feudalism
- |
  feudalist
- |
  feudalistic
- |
  feudalize
- |
  feudally
- |
  feudatory
- |
  fever
- |
  fevered
- |
  feverish
- |
  feverishly
- |
  feverishness
- |
  fewer
- |
  fewness
- |
  feyly
- |
  feyness
- |
  fiance
- |
  fiancee
- |
  fiasco
- |
  fibber
- |
  fiber
- |
  fiberboard
- |
  fiberfill
- |
  Fiberglas
- |
  fiberglass
- |
  fibre
- |
  fibril
- |
  fibrillate
- |
  fibrillation
- |
  fibrin
- |
  fibrinogen
- |
  fibroid
- |
  fibroma
- |
  fibromata
- |
  fibrosis
- |
  fibrotic
- |
  fibrous
- |
  fibula
- |
  fibulae
- |
  fibular
- |
  fiche
- |
  Fichte
- |
  fichu
- |
  fickle
- |
  fickleness
- |
  fickly
- |
  fiction
- |
  fictional
- |
  fictionalize
- |
  fictionally
- |
  fictitious
- |
  fictitiously
- |
  fictive
- |
  fictively
- |
  fictiveness
- |
  ficus
- |
  fiddle
- |
  fiddler
- |
  fiddlestick
- |
  fiddlesticks
- |
  fidelity
- |
  fidget
- |
  fidgetiness
- |
  fidgets
- |
  fidgety
- |
  fiduciary
- |
  Fiedler
- |
  fiefdom
- |
  field
- |
  fielder
- |
  Fielding
- |
  fielding
- |
  Fields
- |
  fieldwork
- |
  fieldworker
- |
  fiend
- |
  fiendish
- |
  fiendishly
- |
  fiendishness
- |
  fierce
- |
  fiercely
- |
  fierceness
- |
  fierily
- |
  fieriness
- |
  fiery
- |
  fiesta
- |
  fifer
- |
  Fifeshire
- |
  fifteen
- |
  fifteenth
- |
  fifth
- |
  fifthly
- |
  fiftieth
- |
  fifty
- |
  Figaro
- |
  fight
- |
  fighter
- |
  fighting
- |
  figment
- |
  figuration
- |
  figurative
- |
  figuratively
- |
  figure
- |
  figurehead
- |
  figurer
- |
  figurine
- |
  Fijian
- |
  filament
- |
  filamentary
- |
  filamented
- |
  filamentous
- |
  filaria
- |
  filariae
- |
  filarial
- |
  filarian
- |
  filbert
- |
  filch
- |
  filcher
- |
  fileable
- |
  filer
- |
  filet
- |
  filial
- |
  filially
- |
  filibuster
- |
  filibusterer
- |
  filigree
- |
  filigreed
- |
  filing
- |
  filings
- |
  Filipino
- |
  filled
- |
  filler
- |
  fillet
- |
  filleter
- |
  filling
- |
  fillip
- |
  Fillmore
- |
  filly
- |
  filmdom
- |
  filmily
- |
  filminess
- |
  filming
- |
  filmmaker
- |
  filmmaking
- |
  filmography
- |
  filmstrip
- |
  filmy
- |
  Filofax
- |
  filter
- |
  filterable
- |
  filterer
- |
  filth
- |
  filthily
- |
  filthiness
- |
  filthy
- |
  filtrable
- |
  filtrate
- |
  filtration
- |
  finagle
- |
  finagler
- |
  final
- |
  finale
- |
  finalise
- |
  finalist
- |
  finality
- |
  finalization
- |
  finalize
- |
  finally
- |
  finance
- |
  finances
- |
  financial
- |
  financially
- |
  financier
- |
  financing
- |
  finch
- |
  findable
- |
  finder
- |
  finding
- |
  finely
- |
  fineness
- |
  finery
- |
  finespun
- |
  finesse
- |
  finfish
- |
  finger
- |
  fingerboard
- |
  fingering
- |
  fingerling
- |
  fingernail
- |
  fingerprint
- |
  fingertip
- |
  finial
- |
  finical
- |
  finickiness
- |
  finicking
- |
  finicky
- |
  finis
- |
  finish
- |
  finished
- |
  finisher
- |
  finite
- |
  finitely
- |
  finiteness
- |
  finitude
- |
  Finland
- |
  Finlander
- |
  finned
- |
  Finnic
- |
  Finnish
- |
  finny
- |
  Fiona
- |
  fiord
- |
  firearm
- |
  fireball
- |
  firebase
- |
  fireboat
- |
  firebomb
- |
  firebox
- |
  firebrand
- |
  firebreak
- |
  firebrick
- |
  firebug
- |
  firecracker
- |
  firedamp
- |
  firedog
- |
  firefight
- |
  firefighter
- |
  firefighting
- |
  firefly
- |
  firehouse
- |
  fireless
- |
  fireman
- |
  Firenze
- |
  fireplace
- |
  fireplug
- |
  firepower
- |
  fireproof
- |
  firer
- |
  fireside
- |
  firestorm
- |
  firetrap
- |
  firetruck
- |
  firewall
- |
  firewater
- |
  firewood
- |
  firework
- |
  fireworks
- |
  firing
- |
  firmament
- |
  firmamental
- |
  firmly
- |
  firmness
- |
  firmware
- |
  first
- |
  firstborn
- |
  firsthand
- |
  firstling
- |
  firstly
- |
  firth
- |
  fiscal
- |
  fiscally
- |
  Fischer
- |
  fishbowl
- |
  fisher
- |
  fisherman
- |
  fishery
- |
  fisheye
- |
  fishhook
- |
  fishily
- |
  fishiness
- |
  fishing
- |
  fishmeal
- |
  fishnet
- |
  fishtail
- |
  fishwife
- |
  fishwives
- |
  fishy
- |
  fissile
- |
  fissility
- |
  fission
- |
  fissionable
- |
  fissure
- |
  fistfight
- |
  fistful
- |
  fisticuff
- |
  fisticuffs
- |
  fistula
- |
  fistulae
- |
  fistulous
- |
  fitful
- |
  fitfully
- |
  fitfulness
- |
  fitly
- |
  fitness
- |
  fitted
- |
  fitter
- |
  fitting
- |
  fittingly
- |
  fittingness
- |
  FitzGerald
- |
  Fitzgerald
- |
  fiver
- |
  fixable
- |
  fixate
- |
  fixated
- |
  fixation
- |
  fixative
- |
  fixed
- |
  fixedly
- |
  fixedness
- |
  fixer
- |
  fixings
- |
  fixity
- |
  fixture
- |
  fizzle
- |
  fizzy
- |
  fjord
- |
  flabbergast
- |
  flabbily
- |
  flabbiness
- |
  flabby
- |
  flaccid
- |
  flaccidity
- |
  flaccidly
- |
  flaccidness
- |
  flack
- |
  flackery
- |
  flacon
- |
  flagella
- |
  flagellar
- |
  flagellate
- |
  flagellation
- |
  flagellator
- |
  flagellatory
- |
  flagellum
- |
  flageolet
- |
  flagger
- |
  flagging
- |
  flagitious
- |
  flagitiously
- |
  flagon
- |
  flagpole
- |
  flagrance
- |
  flagrancy
- |
  flagrant
- |
  flagrantly
- |
  flagship
- |
  flagstaff
- |
  flagstone
- |
  flail
- |
  flair
- |
  flake
- |
  flaker
- |
  flakey
- |
  flakily
- |
  flakiness
- |
  flaky
- |
  flambe
- |
  flambeau
- |
  flambeaux
- |
  flamboyance
- |
  flamboyancy
- |
  flamboyant
- |
  flamboyantly
- |
  flame
- |
  flamenco
- |
  flameout
- |
  flameproof
- |
  flamer
- |
  flamethrower
- |
  flaming
- |
  flamingo
- |
  flammability
- |
  flammable
- |
  Flanders
- |
  flange
- |
  flank
- |
  flanker
- |
  flannel
- |
  flannelet
- |
  flannelette
- |
  flannels
- |
  flapjack
- |
  flapper
- |
  flare
- |
  flareup
- |
  flash
- |
  flashback
- |
  flashbulb
- |
  flashcard
- |
  flashcube
- |
  flasher
- |
  flashgun
- |
  flashily
- |
  flashiness
- |
  flashing
- |
  flashlight
- |
  flashy
- |
  flask
- |
  flatbed
- |
  flatboat
- |
  flatcar
- |
  flatfeet
- |
  flatfish
- |
  flatfoot
- |
  flatfooted
- |
  Flathead
- |
  flatiron
- |
  flatland
- |
  flatly
- |
  flatness
- |
  flats
- |
  flatten
- |
  flattener
- |
  flatter
- |
  flattered
- |
  flatterer
- |
  flattering
- |
  flatteringly
- |
  flattery
- |
  flattish
- |
  flattop
- |
  flatulence
- |
  flatulency
- |
  flatulent
- |
  flatulently
- |
  flatus
- |
  flatware
- |
  flatworm
- |
  Flaubert
- |
  flaunt
- |
  flaunter
- |
  flauntingly
- |
  flaunty
- |
  flautist
- |
  flavor
- |
  flavored
- |
  flavorful
- |
  flavoring
- |
  flavorless
- |
  flavorsome
- |
  flavour
- |
  flavoured
- |
  flawed
- |
  flawless
- |
  flawlessly
- |
  flawlessness
- |
  flaxen
- |
  flayer
- |
  fleabag
- |
  fleabane
- |
  fleck
- |
  flecked
- |
  fledge
- |
  fledgeling
- |
  fledgling
- |
  fleece
- |
  fleeced
- |
  fleecer
- |
  fleecily
- |
  fleeciness
- |
  fleecy
- |
  fleer
- |
  fleeringly
- |
  fleet
- |
  fleeting
- |
  fleetingly
- |
  fleetingness
- |
  fleetly
- |
  fleetness
- |
  Fleming
- |
  Flemish
- |
  flesh
- |
  fleshed
- |
  fleshiness
- |
  fleshliness
- |
  fleshly
- |
  fleshpot
- |
  fleshy
- |
  Fletcher
- |
  flexdollars
- |
  flexibility
- |
  flexible
- |
  flexibleness
- |
  flexibly
- |
  flexitime
- |
  flexor
- |
  flextime
- |
  flexure
- |
  flick
- |
  flicker
- |
  flickeringly
- |
  flied
- |
  flier
- |
  flies
- |
  flight
- |
  flightily
- |
  flightiness
- |
  flightless
- |
  flighty
- |
  flimflam
- |
  flimflammer
- |
  flimflammery
- |
  flimsily
- |
  flimsiness
- |
  flimsy
- |
  flinch
- |
  flincher
- |
  fling
- |
  flinger
- |
  Flint
- |
  flint
- |
  flintily
- |
  flintiness
- |
  flintlock
- |
  flinty
- |
  flippancy
- |
  flippant
- |
  flippantly
- |
  flipper
- |
  flirt
- |
  flirtation
- |
  flirtatious
- |
  flitch
- |
  flitter
- |
  flivver
- |
  float
- |
  floatable
- |
  floater
- |
  floating
- |
  flocculence
- |
  flocculent
- |
  flock
- |
  flocking
- |
  flogger
- |
  flogging
- |
  Flood
- |
  flood
- |
  flooded
- |
  flooder
- |
  floodgate
- |
  flooding
- |
  floodlight
- |
  floodlit
- |
  floodplain
- |
  floodwater
- |
  floor
- |
  floorboard
- |
  flooring
- |
  floorshow
- |
  floorwalker
- |
  floozie
- |
  floozy
- |
  flophouse
- |
  flopper
- |
  floppily
- |
  floppiness
- |
  floppy
- |
  flops
- |
  Flora
- |
  flora
- |
  florae
- |
  floral
- |
  florally
- |
  Florence
- |
  Florentia
- |
  Florentine
- |
  florescence
- |
  florescent
- |
  floret
- |
  florid
- |
  Florida
- |
  Floridan
- |
  Floridian
- |
  floridity
- |
  floridly
- |
  floridness
- |
  florilegia
- |
  florilegium
- |
  florin
- |
  florist
- |
  floruit
- |
  floss
- |
  flossily
- |
  flossiness
- |
  flossy
- |
  flotation
- |
  flotilla
- |
  flotsam
- |
  flounce
- |
  flounced
- |
  flouncy
- |
  flounder
- |
  flour
- |
  flouriness
- |
  flourish
- |
  flourisher
- |
  flourishing
- |
  floury
- |
  flout
- |
  flouter
- |
  flowage
- |
  flowchart
- |
  flower
- |
  flowerbed
- |
  flowered
- |
  flowerily
- |
  floweriness
- |
  flowering
- |
  flowerless
- |
  flowerpot
- |
  flowery
- |
  flowing
- |
  flowingly
- |
  flown
- |
  Floyd
- |
  fluctuant
- |
  fluctuate
- |
  fluctuating
- |
  fluctuation
- |
  fluency
- |
  fluent
- |
  fluently
- |
  fluff
- |
  fluffily
- |
  fluffiness
- |
  fluffy
- |
  fluid
- |
  fluidity
- |
  fluidly
- |
  fluidness
- |
  fluidram
- |
  fluids
- |
  fluke
- |
  flukey
- |
  fluky
- |
  flume
- |
  flummery
- |
  flummox
- |
  flung
- |
  flunk
- |
  flunkey
- |
  flunky
- |
  flunkyism
- |
  fluoresce
- |
  fluorescence
- |
  fluorescent
- |
  fluoridate
- |
  fluoridation
- |
  fluoride
- |
  fluorinate
- |
  fluorination
- |
  fluorine
- |
  fluorite
- |
  fluorocarbon
- |
  fluoroscope
- |
  fluoroscopic
- |
  fluoroscopy
- |
  fluorosis
- |
  flurries
- |
  flurry
- |
  flush
- |
  flushed
- |
  flushness
- |
  fluster
- |
  flustered
- |
  flute
- |
  fluted
- |
  fluting
- |
  flutist
- |
  flutter
- |
  fluttery
- |
  fluty
- |
  fluvial
- |
  flyable
- |
  flyblown
- |
  flyby
- |
  flycatcher
- |
  flyer
- |
  flying
- |
  flyleaf
- |
  flyleaves
- |
  flypaper
- |
  flyspeck
- |
  flyswatter
- |
  flyway
- |
  flyweight
- |
  flywheel
- |
  foaminess
- |
  foamy
- |
  focaccia
- |
  focal
- |
  focally
- |
  focus
- |
  fodder
- |
  foehn
- |
  foeman
- |
  foetal
- |
  foetid
- |
  foetus
- |
  fogbound
- |
  fogey
- |
  fogeydom
- |
  fogeyish
- |
  fogeyism
- |
  foggily
- |
  fogginess
- |
  foggy
- |
  foghorn
- |
  fogyish
- |
  foible
- |
  foilist
- |
  foist
- |
  Fokine
- |
  foldable
- |
  foldaway
- |
  folder
- |
  folderol
- |
  foldout
- |
  foliage
- |
  foliate
- |
  foliated
- |
  folio
- |
  folklore
- |
  folkloric
- |
  folklorist
- |
  folkloristic
- |
  folks
- |
  folksiness
- |
  folksinger
- |
  folksinging
- |
  folksong
- |
  folksy
- |
  folkway
- |
  follicle
- |
  follies
- |
  follow
- |
  follower
- |
  following
- |
  followup
- |
  folly
- |
  Fomalhaut
- |
  foment
- |
  fomentation
- |
  fomenter
- |
  Fonda
- |
  fondant
- |
  fondle
- |
  fondly
- |
  fondness
- |
  fondu
- |
  fondue
- |
  fontanel
- |
  fontanelle
- |
  Fonteyn
- |
  Foochow
- |
  foodie
- |
  foodstuff
- |
  foolery
- |
  foolhardily
- |
  foolhardy
- |
  foolish
- |
  foolishly
- |
  foolishness
- |
  foolproof
- |
  foolscap
- |
  footage
- |
  football
- |
  footballer
- |
  footballing
- |
  footboard
- |
  footbridge
- |
  footed
- |
  footfall
- |
  footgear
- |
  foothill
- |
  foothills
- |
  foothold
- |
  footing
- |
  footless
- |
  footlessly
- |
  footlessness
- |
  footlights
- |
  footling
- |
  footlocker
- |
  footloose
- |
  footman
- |
  footnote
- |
  footpad
- |
  footpath
- |
  footprint
- |
  footrace
- |
  footrest
- |
  footsie
- |
  footsore
- |
  footsoreness
- |
  footstep
- |
  footstool
- |
  footwear
- |
  footwork
- |
  foppery
- |
  foppish
- |
  foppishly
- |
  foppishness
- |
  forage
- |
  forager
- |
  Foraker
- |
  foray
- |
  forayer
- |
  forbad
- |
  forbade
- |
  forbear
- |
  forbearance
- |
  forbearer
- |
  forbid
- |
  forbiddance
- |
  forbidden
- |
  forbidding
- |
  forbiddingly
- |
  forbode
- |
  forbore
- |
  forborne
- |
  force
- |
  forced
- |
  forcedly
- |
  forceful
- |
  forcefully
- |
  forcefulness
- |
  forceless
- |
  forceps
- |
  forcer
- |
  forces
- |
  forcible
- |
  forcibly
- |
  fordable
- |
  forearm
- |
  forebear
- |
  forebode
- |
  foreboding
- |
  forebodingly
- |
  forecast
- |
  forecaster
- |
  forecastle
- |
  foreclose
- |
  foreclosure
- |
  forecourt
- |
  foredoom
- |
  forefather
- |
  forefathers
- |
  forefeet
- |
  forefend
- |
  forefinger
- |
  forefoot
- |
  forefront
- |
  foregather
- |
  forego
- |
  foregoer
- |
  foregoing
- |
  foregone
- |
  foreground
- |
  forehand
- |
  forehanded
- |
  forehead
- |
  foreign
- |
  foreigner
- |
  foreignness
- |
  foreknew
- |
  foreknow
- |
  foreknown
- |
  forelady
- |
  foreleg
- |
  forelimb
- |
  forelock
- |
  foreman
- |
  foremast
- |
  foremost
- |
  forename
- |
  forenamed
- |
  forenoon
- |
  forensic
- |
  forensically
- |
  forensics
- |
  foreordain
- |
  forepart
- |
  foreperson
- |
  foreplay
- |
  forequarter
- |
  forerunner
- |
  foresail
- |
  foresaw
- |
  foresee
- |
  foreseeable
- |
  foreseen
- |
  foreseer
- |
  foreshadow
- |
  foreshadower
- |
  foreshore
- |
  foreshorten
- |
  foresight
- |
  foresighted
- |
  foreskin
- |
  Forest
- |
  forest
- |
  forestall
- |
  forestation
- |
  forested
- |
  forester
- |
  forestland
- |
  forestry
- |
  foreswear
- |
  foretaste
- |
  foretell
- |
  foreteller
- |
  forethought
- |
  foretoken
- |
  foretold
- |
  foretop
- |
  forever
- |
  forevermore
- |
  forewarn
- |
  forewent
- |
  forewing
- |
  forewoman
- |
  foreword
- |
  forfeit
- |
  forfeitable
- |
  forfeiter
- |
  forfeiture
- |
  forfend
- |
  forgather
- |
  forgave
- |
  forge
- |
  forger
- |
  forgery
- |
  forget
- |
  forgetful
- |
  forgetfully
- |
  forgettable
- |
  forging
- |
  forgivable
- |
  forgive
- |
  forgiven
- |
  forgiveness
- |
  forgiver
- |
  forgiving
- |
  forgivingly
- |
  forgo
- |
  forgoer
- |
  forgone
- |
  forgot
- |
  forgotten
- |
  forint
- |
  forked
- |
  forkful
- |
  forklift
- |
  forlorn
- |
  forlornly
- |
  forlornness
- |
  formal
- |
  formaldehyde
- |
  formalise
- |
  formalism
- |
  formalist
- |
  formalistic
- |
  formalities
- |
  formality
- |
  formalize
- |
  formally
- |
  format
- |
  formation
- |
  formational
- |
  formative
- |
  formatted
- |
  formatter
- |
  formatting
- |
  former
- |
  formerly
- |
  formfitting
- |
  formic
- |
  Formica
- |
  formication
- |
  formidable
- |
  formidably
- |
  formless
- |
  formlessly
- |
  formlessness
- |
  Formosa
- |
  Formosan
- |
  formula
- |
  formulae
- |
  formulaic
- |
  formulate
- |
  formulation
- |
  formulator
- |
  Fornax
- |
  fornicate
- |
  fornication
- |
  fornicator
- |
  Forrest
- |
  forsake
- |
  forsaken
- |
  forsook
- |
  forsooth
- |
  Forster
- |
  forswear
- |
  forswore
- |
  forsworn
- |
  Forsyth
- |
  forsythia
- |
  Fortaleza
- |
  forte
- |
  Forth
- |
  forth
- |
  forthcoming
- |
  forthright
- |
  forthrightly
- |
  forthwith
- |
  fortieth
- |
  fortified
- |
  fortifier
- |
  fortify
- |
  fortissimo
- |
  fortitude
- |
  fortnight
- |
  fortnightly
- |
  FORTRAN
- |
  fortress
- |
  fortuitous
- |
  fortuitously
- |
  fortuity
- |
  fortunate
- |
  fortunately
- |
  fortune
- |
  fortunes
- |
  forty
- |
  forum
- |
  forward
- |
  forwarder
- |
  forwarding
- |
  forwardly
- |
  forwardness
- |
  forwards
- |
  forwent
- |
  fossil
- |
  fossilize
- |
  Foster
- |
  foster
- |
  fosterling
- |
  Foucault
- |
  fought
- |
  foulard
- |
  foully
- |
  foulmouthed
- |
  foulness
- |
  found
- |
  foundation
- |
  foundational
- |
  founded
- |
  founder
- |
  founding
- |
  foundling
- |
  foundry
- |
  fount
- |
  fountain
- |
  fountainhead
- |
  fourfold
- |
  Fourier
- |
  fourposter
- |
  fourscore
- |
  foursome
- |
  foursquare
- |
  fourteen
- |
  fourteenth
- |
  fourth
- |
  fourthly
- |
  fourwheeled
- |
  Fowles
- |
  foxed
- |
  foxfire
- |
  foxglove
- |
  foxhole
- |
  foxhound
- |
  foxily
- |
  foxiness
- |
  foxtrot
- |
  foyer
- |
  frabjous
- |
  fracas
- |
  fractal
- |
  fraction
- |
  fractional
- |
  fractionally
- |
  fractious
- |
  fractiously
- |
  fracture
- |
  fractured
- |
  fragile
- |
  fragilely
- |
  fragileness
- |
  fragility
- |
  fragment
- |
  fragmental
- |
  fragmentary
- |
  fragmented
- |
  Fragonard
- |
  fragrance
- |
  fragrant
- |
  fragrantly
- |
  frail
- |
  frailly
- |
  frailness
- |
  frailty
- |
  frame
- |
  framer
- |
  frames
- |
  framework
- |
  franc
- |
  France
- |
  Frances
- |
  franchisable
- |
  franchise
- |
  franchisee
- |
  franchiser
- |
  franchising
- |
  franchisor
- |
  Francine
- |
  Francis
- |
  Franciscan
- |
  Francisco
- |
  francium
- |
  Franck
- |
  Franco
- |
  Francophone
- |
  francophone
- |
  frangibility
- |
  frangible
- |
  Frank
- |
  frank
- |
  Frankenstein
- |
  Frankfort
- |
  Frankfurt
- |
  frankfurt
- |
  Frankfurter
- |
  frankfurter
- |
  frankincense
- |
  Frankish
- |
  Franklin
- |
  frankly
- |
  Franklyn
- |
  frankness
- |
  frantic
- |
  frantically
- |
  franticly
- |
  frappe
- |
  Fraser
- |
  fraternal
- |
  fraternalism
- |
  fraternally
- |
  fraternity
- |
  fraternize
- |
  fraternizer
- |
  fratricidal
- |
  fratricide
- |
  fraud
- |
  fraudulence
- |
  fraudulent
- |
  fraudulently
- |
  Frauen
- |
  fraught
- |
  Fraulein
- |
  frayed
- |
  Frazer
- |
  frazzle
- |
  frazzled
- |
  freak
- |
  freakily
- |
  freakish
- |
  freakishly
- |
  freakishness
- |
  freakout
- |
  freaky
- |
  freckle
- |
  freckled
- |
  freckly
- |
  Freda
- |
  Freddie
- |
  Frederic
- |
  Frederica
- |
  Frederick
- |
  Fredericka
- |
  Fredericton
- |
  Fredric
- |
  Fredrick
- |
  freebase
- |
  freebee
- |
  freebie
- |
  freeboard
- |
  freeboot
- |
  freebooter
- |
  freeborn
- |
  freedman
- |
  freedom
- |
  freedwoman
- |
  freeform
- |
  freehand
- |
  freehanded
- |
  freehandedly
- |
  freehold
- |
  freeholder
- |
  freelance
- |
  freelancer
- |
  freeload
- |
  freeloader
- |
  freely
- |
  Freeman
- |
  freeman
- |
  Freemason
- |
  Freemasonry
- |
  freeness
- |
  freestanding
- |
  freestone
- |
  freestyle
- |
  freethinker
- |
  freethinking
- |
  Freetown
- |
  freeware
- |
  freeway
- |
  freewheel
- |
  freewheeling
- |
  freewill
- |
  freezable
- |
  freeze
- |
  freezer
- |
  freezing
- |
  freight
- |
  freighter
- |
  Fremont
- |
  frena
- |
  French
- |
  Frenchman
- |
  Frenchwoman
- |
  frenetic
- |
  frenetical
- |
  frenetically
- |
  frenum
- |
  frenzied
- |
  frenziedly
- |
  frenzy
- |
  Freon
- |
  frequency
- |
  frequent
- |
  frequenter
- |
  frequently
- |
  frequentness
- |
  fresco
- |
  fresh
- |
  freshen
- |
  freshener
- |
  freshet
- |
  freshly
- |
  freshman
- |
  freshness
- |
  freshwater
- |
  Fresno
- |
  fretful
- |
  fretfully
- |
  fretfulness
- |
  fretsaw
- |
  fretted
- |
  fretter
- |
  fretwork
- |
  Freud
- |
  Freudian
- |
  Freudianism
- |
  Freya
- |
  Freyja
- |
  Freyr
- |
  friability
- |
  friable
- |
  friableness
- |
  friar
- |
  friary
- |
  fricassee
- |
  fricative
- |
  friction
- |
  frictional
- |
  frictionally
- |
  frictionless
- |
  Friday
- |
  fridge
- |
  fried
- |
  Frieda
- |
  Friedan
- |
  friedcake
- |
  Friedman
- |
  Friend
- |
  friend
- |
  friendless
- |
  friendlily
- |
  friendliness
- |
  friendly
- |
  friendship
- |
  frier
- |
  fries
- |
  frieze
- |
  frigate
- |
  Frigga
- |
  frigging
- |
  fright
- |
  frighten
- |
  frightened
- |
  frightening
- |
  frightful
- |
  frightfully
- |
  frigid
- |
  frigidity
- |
  frigidly
- |
  frigidness
- |
  frill
- |
  frilliness
- |
  frilly
- |
  Friml
- |
  fringe
- |
  fringed
- |
  fringy
- |
  frippery
- |
  Frisbee
- |
  frise
- |
  Frisian
- |
  frisk
- |
  frisker
- |
  friskily
- |
  friskiness
- |
  frisky
- |
  frisson
- |
  frittata
- |
  fritter
- |
  Fritz
- |
  fritz
- |
  frivolity
- |
  frivolous
- |
  frivolously
- |
  frizz
- |
  frizzle
- |
  frizzly
- |
  frizzy
- |
  Frobisher
- |
  frock
- |
  frogman
- |
  froideur
- |
  Froissart
- |
  frolic
- |
  frolicker
- |
  frolicsome
- |
  frond
- |
  front
- |
  frontage
- |
  frontal
- |
  frontally
- |
  Frontenac
- |
  frontier
- |
  frontiersman
- |
  frontispiece
- |
  frontline
- |
  frontrunner
- |
  frontward
- |
  frontwards
- |
  frosh
- |
  Frost
- |
  frost
- |
  frostbit
- |
  frostbite
- |
  frostbitten
- |
  frostily
- |
  frostiness
- |
  frosting
- |
  frosty
- |
  froth
- |
  frothily
- |
  frothiness
- |
  frothy
- |
  frottage
- |
  frotteur
- |
  frotteurism
- |
  froufrou
- |
  Froward
- |
  froward
- |
  frowardly
- |
  frowardness
- |
  frown
- |
  frowner
- |
  frowningly
- |
  frowsy
- |
  frowzily
- |
  frowziness
- |
  frowzy
- |
  froze
- |
  frozen
- |
  fructiferous
- |
  fructify
- |
  fructose
- |
  fructuous
- |
  frugal
- |
  frugality
- |
  frugally
- |
  frugalness
- |
  fruit
- |
  fruitarian
- |
  fruitcake
- |
  fruited
- |
  fruitful
- |
  fruitfully
- |
  fruitfulness
- |
  fruitily
- |
  fruitiness
- |
  fruition
- |
  fruitless
- |
  fruitlessly
- |
  fruity
- |
  frump
- |
  frumpily
- |
  frumpiness
- |
  frumpish
- |
  frumpishly
- |
  frumpishness
- |
  frumpy
- |
  Frunze
- |
  frusta
- |
  frustrate
- |
  frustrated
- |
  frustrater
- |
  frustrating
- |
  frustration
- |
  frustum
- |
  fryable
- |
  fryer
- |
  Fuchou
- |
  fuchsia
- |
  fucker
- |
  fucking
- |
  fuddle
- |
  fudge
- |
  fuehrer
- |
  fueler
- |
  Fuentes
- |
  fugacious
- |
  fugaciously
- |
  fugal
- |
  fugally
- |
  fugitive
- |
  fugue
- |
  fuguist
- |
  Fuhrer
- |
  fuhrer
- |
  Fujiyama
- |
  Fukuoka
- |
  Fulbright
- |
  fulcra
- |
  fulcrum
- |
  fulfil
- |
  fulfill
- |
  fulfilled
- |
  fulfiller
- |
  fulfilling
- |
  fulfillment
- |
  fulfilment
- |
  fulgurant
- |
  fulgurate
- |
  fulguration
- |
  fulgurous
- |
  fuliginous
- |
  fullback
- |
  Fuller
- |
  fuller
- |
  fullerene
- |
  Fullerton
- |
  fulling
- |
  fullness
- |
  fully
- |
  fulminant
- |
  fulminate
- |
  fulminating
- |
  fulmination
- |
  fulminator
- |
  fulminatory
- |
  fulness
- |
  fulsome
- |
  fulsomely
- |
  fulsomeness
- |
  Fulton
- |
  fulvous
- |
  fumarole
- |
  fumble
- |
  fumbler
- |
  fumblingly
- |
  fumes
- |
  fumigant
- |
  fumigate
- |
  fumigation
- |
  fumigator
- |
  Funabashi
- |
  Funafuti
- |
  funambulist
- |
  function
- |
  functional
- |
  functionally
- |
  functionary
- |
  functionless
- |
  fundament
- |
  fundamental
- |
  fundamentals
- |
  funding
- |
  fundraiser
- |
  fundraising
- |
  funds
- |
  Fundy
- |
  funeral
- |
  funerary
- |
  funereal
- |
  funereally
- |
  fungal
- |
  fungi
- |
  fungibility
- |
  fungible
- |
  fungicidal
- |
  fungicide
- |
  fungo
- |
  fungous
- |
  fungus
- |
  funicular
- |
  funkily
- |
  funkiness
- |
  funky
- |
  funnel
- |
  funnies
- |
  funnily
- |
  funniness
- |
  funny
- |
  furbelow
- |
  furbelowed
- |
  furbelows
- |
  furbish
- |
  Furies
- |
  furious
- |
  furiously
- |
  furlong
- |
  furlough
- |
  furnace
- |
  furnish
- |
  furnished
- |
  furnisher
- |
  furnishings
- |
  furniture
- |
  furor
- |
  furore
- |
  furred
- |
  furrier
- |
  furriness
- |
  furring
- |
  furrow
- |
  furrowed
- |
  furry
- |
  further
- |
  furtherance
- |
  furthermore
- |
  furthermost
- |
  furthest
- |
  furtive
- |
  furtively
- |
  furtiveness
- |
  furze
- |
  furzy
- |
  fuscous
- |
  fusebox
- |
  fusee
- |
  fuselage
- |
  Fushun
- |
  fusibility
- |
  fusible
- |
  fusileer
- |
  fusilier
- |
  fusillade
- |
  fusion
- |
  fusional
- |
  fussbudget
- |
  fusser
- |
  fussily
- |
  fussiness
- |
  fusspot
- |
  fussy
- |
  fustian
- |
  fustily
- |
  fustiness
- |
  fusty
- |
  futile
- |
  futilely
- |
  futility
- |
  futon
- |
  future
- |
  futures
- |
  Futurism
- |
  futurism
- |
  futurist
- |
  futuristic
- |
  futurity
- |
  futurologist
- |
  futurology
- |
  fuzee
- |
  Fuzhou
- |
  fuzzily
- |
  fuzziness
- |
  fuzzy
- |
  gabardine
- |
  gabber
- |
  gabbiness
- |
  gabble
- |
  gabbler
- |
  gabby
- |
  gaberdine
- |
  gabfest
- |
  Gable
- |
  gable
- |
  gabled
- |
  Gabon
- |
  Gabonese
- |
  Gaborone
- |
  Gabriel
- |
  Gabrielle
- |
  gadabout
- |
  Gaddafi
- |
  gadder
- |
  gadfly
- |
  gadget
- |
  gadgetry
- |
  gadolinium
- |
  Gaelic
- |
  gaffe
- |
  gaffer
- |
  Gagarin
- |
  gagged
- |
  gagger
- |
  gaggle
- |
  gaiety
- |
  gaily
- |
  gainer
- |
  Gainesville
- |
  gainful
- |
  gainfully
- |
  gains
- |
  gainsaid
- |
  gainsay
- |
  gainsayer
- |
  Gainsborough
- |
  gaited
- |
  gaiter
- |
  galabia
- |
  galabiya
- |
  galactic
- |
  galactose
- |
  Galahad
- |
  Galatea
- |
  Galatia
- |
  Galatian
- |
  Galatians
- |
  Galaxy
- |
  galaxy
- |
  Galbraith
- |
  Galen
- |
  galena
- |
  galere
- |
  Galicia
- |
  Galician
- |
  Galilean
- |
  Galilee
- |
  Galilei
- |
  Galileo
- |
  gallant
- |
  gallantly
- |
  gallantries
- |
  gallantry
- |
  gallbladder
- |
  galleon
- |
  galleria
- |
  galleried
- |
  gallery
- |
  galley
- |
  galliard
- |
  Gallic
- |
  Gallicism
- |
  gallimaufry
- |
  galling
- |
  gallinule
- |
  gallium
- |
  gallivant
- |
  gallon
- |
  gallop
- |
  galloper
- |
  galloping
- |
  Galloway
- |
  gallows
- |
  gallstone
- |
  Gallup
- |
  galluses
- |
  galore
- |
  galosh
- |
  galoshe
- |
  galoshes
- |
  Galsworthy
- |
  galumph
- |
  Galvani
- |
  galvanic
- |
  galvanically
- |
  galvanise
- |
  galvanism
- |
  galvanize
- |
  galvanized
- |
  galvanizer
- |
  galvanometer
- |
  Galveston
- |
  Galway
- |
  gambade
- |
  gambado
- |
  Gambia
- |
  Gambian
- |
  gambit
- |
  gamble
- |
  gambler
- |
  gambling
- |
  gambol
- |
  gambrel
- |
  gamecock
- |
  gamekeeper
- |
  gamely
- |
  gameness
- |
  games
- |
  gamesmanship
- |
  gamesome
- |
  gamester
- |
  gamete
- |
  gametic
- |
  gamey
- |
  gamin
- |
  gamine
- |
  gaminess
- |
  gaming
- |
  gamma
- |
  gammer
- |
  gammon
- |
  gamut
- |
  gander
- |
  Gandhi
- |
  gangbusters
- |
  Ganges
- |
  Gangetic
- |
  gangland
- |
  ganglia
- |
  gangling
- |
  ganglion
- |
  ganglionic
- |
  gangly
- |
  gangplank
- |
  gangplow
- |
  gangrene
- |
  gangrenous
- |
  gangster
- |
  gangsterdom
- |
  gangsterism
- |
  gangway
- |
  ganja
- |
  gannet
- |
  gantlet
- |
  gantry
- |
  gaoler
- |
  gaping
- |
  gappy
- |
  garage
- |
  garbage
- |
  garbageman
- |
  garbanzo
- |
  garble
- |
  garbled
- |
  garbler
- |
  Garbo
- |
  garbologist
- |
  garbology
- |
  garcon
- |
  garden
- |
  gardener
- |
  gardenia
- |
  gardening
- |
  gardens
- |
  garderobe
- |
  Gardner
- |
  Garfield
- |
  garfish
- |
  Gargantua
- |
  Gargantuan
- |
  gargantuan
- |
  gargle
- |
  gargoyle
- |
  gargoyled
- |
  Garibaldi
- |
  garish
- |
  garishly
- |
  garishness
- |
  Garland
- |
  garland
- |
  garlic
- |
  garlicky
- |
  garment
- |
  garner
- |
  garnet
- |
  garnish
- |
  garnishee
- |
  garnishment
- |
  garniture
- |
  Garonne
- |
  garote
- |
  garotte
- |
  garret
- |
  Garrett
- |
  Garrick
- |
  Garrison
- |
  garrison
- |
  garrote
- |
  garroter
- |
  garrotte
- |
  garrulity
- |
  garrulous
- |
  garrulously
- |
  Garry
- |
  garter
- |
  Garth
- |
  Garvey
- |
  Gascon
- |
  gasconade
- |
  Gascony
- |
  gaseous
- |
  gasket
- |
  gaslight
- |
  gasohol
- |
  gasolene
- |
  gasoline
- |
  Gaspe
- |
  Gaspesian
- |
  gassiness
- |
  gassy
- |
  gastric
- |
  gastritis
- |
  gastrologic
- |
  gastrologist
- |
  gastrology
- |
  gastronome
- |
  gastronomic
- |
  gastronomy
- |
  gastropod
- |
  gasworks
- |
  gatecrash
- |
  gatecrasher
- |
  gated
- |
  gatefold
- |
  gatehouse
- |
  gatekeeper
- |
  gatepost
- |
  gater
- |
  Gates
- |
  Gateshead
- |
  gateway
- |
  gather
- |
  gathered
- |
  gatherer
- |
  gathering
- |
  gathers
- |
  gator
- |
  gauche
- |
  gauchely
- |
  gaucheness
- |
  gaucherie
- |
  gaucho
- |
  gaudily
- |
  gaudiness
- |
  gaudy
- |
  gauge
- |
  gaugeable
- |
  gauged
- |
  gauger
- |
  Gauguin
- |
  Gauhati
- |
  Gaulish
- |
  Gaullism
- |
  Gaullist
- |
  gaunt
- |
  gauntlet
- |
  gauntly
- |
  gauntness
- |
  Gautama
- |
  Gautier
- |
  gauze
- |
  gauzily
- |
  gauziness
- |
  gauzy
- |
  gavage
- |
  gavel
- |
  gavotte
- |
  Gawain
- |
  gawker
- |
  gawkily
- |
  gawkiness
- |
  gawky
- |
  gayety
- |
  Gayle
- |
  Gaylord
- |
  gayly
- |
  gayness
- |
  gazebo
- |
  gazelle
- |
  gazer
- |
  gazette
- |
  gazetteer
- |
  Gaziantep
- |
  gazpacho
- |
  Gdansk
- |
  Gdynia
- |
  gearbox
- |
  gearshift
- |
  gearwheel
- |
  gecko
- |
  geegaw
- |
  geeky
- |
  Geelong
- |
  geese
- |
  geezer
- |
  gegenschein
- |
  Gehrig
- |
  geisha
- |
  gelatin
- |
  gelatine
- |
  gelatinous
- |
  gelcap
- |
  gelding
- |
  gelid
- |
  gelidity
- |
  gelidness
- |
  gelignite
- |
  geminate
- |
  geminately
- |
  gemination
- |
  Gemini
- |
  gemmologist
- |
  gemmology
- |
  gemmy
- |
  gemological
- |
  gemologist
- |
  gemology
- |
  gemstone
- |
  gemutlich
- |
  gendarme
- |
  gendarmerie
- |
  gender
- |
  genderless
- |
  genealogical
- |
  genealogist
- |
  genealogize
- |
  genealogy
- |
  genera
- |
  general
- |
  generalise
- |
  generalised
- |
  generalist
- |
  generality
- |
  generalize
- |
  generalized
- |
  generally
- |
  generalship
- |
  generate
- |
  generation
- |
  generational
- |
  generative
- |
  generator
- |
  generic
- |
  generically
- |
  generosity
- |
  generous
- |
  generously
- |
  generousness
- |
  geneses
- |
  Genesis
- |
  genesis
- |
  Genet
- |
  genetic
- |
  genetically
- |
  geneticist
- |
  genetics
- |
  Geneva
- |
  Genevan
- |
  Genevese
- |
  Genevieve
- |
  Genghis
- |
  genial
- |
  geniality
- |
  genially
- |
  genialness
- |
  genic
- |
  genie
- |
  genii
- |
  genital
- |
  genitalia
- |
  genitalic
- |
  genitally
- |
  genitals
- |
  genitival
- |
  genitivally
- |
  genitive
- |
  genius
- |
  Genoa
- |
  genocidal
- |
  genocidally
- |
  genocide
- |
  Genoese
- |
  genome
- |
  genomic
- |
  genomics
- |
  genotype
- |
  genotypic
- |
  genotypical
- |
  Genovese
- |
  genre
- |
  genteel
- |
  genteelly
- |
  genteelness
- |
  gentes
- |
  gentian
- |
  Gentile
- |
  gentile
- |
  gentility
- |
  gentle
- |
  gentlefolk
- |
  gentlefolks
- |
  gentleman
- |
  gentlemanly
- |
  gentleness
- |
  gentlewoman
- |
  gently
- |
  gentrified
- |
  gentrifier
- |
  gentrify
- |
  gentry
- |
  genuflect
- |
  genuflection
- |
  genuflector
- |
  genuflexion
- |
  genuine
- |
  genuinely
- |
  genuineness
- |
  genus
- |
  geocentric
- |
  geocentrism
- |
  geochemical
- |
  geochemist
- |
  geochemistry
- |
  geode
- |
  geodesic
- |
  geodesist
- |
  geodesy
- |
  geodetic
- |
  Geoffrey
- |
  geographer
- |
  geographic
- |
  geographical
- |
  geography
- |
  geologic
- |
  geological
- |
  geologically
- |
  geologist
- |
  geology
- |
  geomagnetic
- |
  geomagnetism
- |
  geomancer
- |
  geomancy
- |
  geomantic
- |
  geometer
- |
  Geometric
- |
  geometric
- |
  geometrical
- |
  geometrician
- |
  geometry
- |
  geophysical
- |
  geophysicist
- |
  geophysics
- |
  geopolitical
- |
  geopolitics
- |
  George
- |
  Georgeann
- |
  Georgetown
- |
  Georgette
- |
  Georgia
- |
  Georgian
- |
  georgic
- |
  Georgics
- |
  Georgina
- |
  geosyncline
- |
  geothermal
- |
  geothermally
- |
  geothermic
- |
  Gerald
- |
  Geraldine
- |
  geranium
- |
  Gerard
- |
  gerbil
- |
  gerbile
- |
  Gerhard
- |
  geriatric
- |
  geriatrics
- |
  German
- |
  germane
- |
  germanely
- |
  germaneness
- |
  Germanic
- |
  germanium
- |
  Germantown
- |
  Germany
- |
  germicidal
- |
  germicide
- |
  germinable
- |
  germinal
- |
  germinally
- |
  germinate
- |
  germination
- |
  germinative
- |
  germinator
- |
  germy
- |
  Geronimo
- |
  gerontocracy
- |
  gerontocrat
- |
  gerontologic
- |
  gerontology
- |
  Gerry
- |
  gerrymander
- |
  Gershwin
- |
  Gertrude
- |
  gerund
- |
  gerundial
- |
  gerundive
- |
  Gestalt
- |
  gestalt
- |
  Gestalten
- |
  gestalten
- |
  gestaltism
- |
  gestaltist
- |
  Gestapo
- |
  gestapo
- |
  gestate
- |
  gestation
- |
  gestational
- |
  gestatory
- |
  gesticulate
- |
  gesticulator
- |
  gestural
- |
  gesture
- |
  gesturer
- |
  gesundheit
- |
  getaway
- |
  Getty
- |
  Gettysburg
- |
  getup
- |
  gewgaw
- |
  geyser
- |
  Ghana
- |
  Ghanaian
- |
  Ghanian
- |
  ghastliness
- |
  ghastly
- |
  Ghats
- |
  Ghent
- |
  gherkin
- |
  ghetto
- |
  ghettoize
- |
  ghost
- |
  ghostliness
- |
  ghostly
- |
  ghostwrite
- |
  ghostwriter
- |
  ghostwriting
- |
  ghostwritten
- |
  ghostwrote
- |
  ghoul
- |
  ghoulish
- |
  ghoulishly
- |
  ghoulishness
- |
  Giacometti
- |
  giant
- |
  giantess
- |
  gibber
- |
  gibbering
- |
  gibberish
- |
  gibbet
- |
  Gibbon
- |
  gibbon
- |
  gibbosity
- |
  gibbous
- |
  gibbously
- |
  gibbousness
- |
  giber
- |
  gibingly
- |
  giblet
- |
  giblets
- |
  Gibraltar
- |
  Gibson
- |
  giddily
- |
  giddiness
- |
  giddy
- |
  Gideon
- |
  Gielgud
- |
  gifted
- |
  giftedness
- |
  gigabyte
- |
  gigaflops
- |
  gigahertz
- |
  gigantic
- |
  gigantically
- |
  gigantism
- |
  giggle
- |
  giggler
- |
  giggly
- |
  gigolo
- |
  Gijon
- |
  Gilbert
- |
  Gilda
- |
  gilder
- |
  gilding
- |
  Gilead
- |
  Gileadite
- |
  Giles
- |
  gilled
- |
  Gillespie
- |
  Gillian
- |
  gillyflower
- |
  Gilman
- |
  gimbal
- |
  gimbals
- |
  gimcrack
- |
  gimcrackery
- |
  gimlet
- |
  gimme
- |
  gimmick
- |
  gimmickry
- |
  gimmicky
- |
  gimpy
- |
  Ginger
- |
  ginger
- |
  gingerbread
- |
  gingerliness
- |
  gingerly
- |
  gingersnap
- |
  gingery
- |
  gingham
- |
  gingiva
- |
  gingivae
- |
  gingivitis
- |
  gingko
- |
  ginkgo
- |
  ginny
- |
  Ginsberg
- |
  Ginsburg
- |
  ginseng
- |
  Giorgione
- |
  Giotto
- |
  Gipsy
- |
  gipsy
- |
  giraffe
- |
  Giraudoux
- |
  girder
- |
  girdle
- |
  girdler
- |
  girlfriend
- |
  girlhood
- |
  girlish
- |
  girlishly
- |
  girlishness
- |
  girly
- |
  girth
- |
  Gisela
- |
  Giselle
- |
  gismo
- |
  giveaway
- |
  giveback
- |
  given
- |
  giver
- |
  giving
- |
  gizmo
- |
  gizzard
- |
  glabrous
- |
  glace
- |
  glacial
- |
  glacially
- |
  glaciate
- |
  glaciation
- |
  glacier
- |
  glacis
- |
  gladden
- |
  glade
- |
  gladiator
- |
  gladiatorial
- |
  gladiola
- |
  gladioli
- |
  gladiolus
- |
  gladly
- |
  gladness
- |
  gladsome
- |
  gladsomely
- |
  Gladstone
- |
  gladstone
- |
  Gladys
- |
  glamor
- |
  glamorize
- |
  glamorizer
- |
  glamorous
- |
  glamorously
- |
  glamour
- |
  glamourize
- |
  glamourous
- |
  glance
- |
  glancing
- |
  glancingly
- |
  gland
- |
  glandes
- |
  glandular
- |
  glandularly
- |
  glans
- |
  glare
- |
  glaring
- |
  glaringly
- |
  Glasgow
- |
  glasnost
- |
  glass
- |
  glassblower
- |
  glassblowing
- |
  glasses
- |
  glassful
- |
  glassily
- |
  glassiness
- |
  glassware
- |
  glassy
- |
  Glaswegian
- |
  glaucoma
- |
  glaucous
- |
  glaze
- |
  glazed
- |
  glazer
- |
  glazier
- |
  glaziery
- |
  gleam
- |
  gleamy
- |
  glean
- |
  gleanable
- |
  gleaner
- |
  gleaning
- |
  gleanings
- |
  Gleason
- |
  gleeful
- |
  gleefully
- |
  gleefulness
- |
  Glenda
- |
  Glendale
- |
  Glendower
- |
  glengarry
- |
  Glenn
- |
  Glenna
- |
  glibly
- |
  glibness
- |
  glide
- |
  glider
- |
  gliding
- |
  glimmer
- |
  glimmering
- |
  glimpse
- |
  glint
- |
  glissade
- |
  glissandi
- |
  glissando
- |
  glisten
- |
  glistening
- |
  glister
- |
  glitch
- |
  glitchy
- |
  glitter
- |
  glitterati
- |
  glittering
- |
  glitteringly
- |
  glittery
- |
  glitz
- |
  glitzily
- |
  glitziness
- |
  glitzy
- |
  gloaming
- |
  gloat
- |
  gloater
- |
  gloatingly
- |
  global
- |
  globalism
- |
  globalist
- |
  globalize
- |
  globally
- |
  globe
- |
  globetrot
- |
  globetrotter
- |
  globular
- |
  globularly
- |
  globularness
- |
  globule
- |
  globulin
- |
  globulous
- |
  glockenspiel
- |
  gloom
- |
  gloomily
- |
  gloominess
- |
  gloomy
- |
  gloppy
- |
  Gloria
- |
  glorified
- |
  glorifier
- |
  glorify
- |
  glorious
- |
  gloriously
- |
  gloriousness
- |
  glory
- |
  gloss
- |
  glossarial
- |
  glossary
- |
  glosser
- |
  glossily
- |
  glossiness
- |
  glossolalia
- |
  glossolalic
- |
  glossy
- |
  glottal
- |
  glottides
- |
  glottis
- |
  Gloucester
- |
  glove
- |
  glower
- |
  glowering
- |
  gloweringly
- |
  glowing
- |
  glowingly
- |
  glowworm
- |
  gloxinia
- |
  gloze
- |
  glucagon
- |
  glucose
- |
  gluey
- |
  gluiness
- |
  glumly
- |
  glumness
- |
  gluon
- |
  gluteal
- |
  glutei
- |
  gluten
- |
  glutenous
- |
  gluteus
- |
  glutinosity
- |
  glutinous
- |
  glutinously
- |
  glutton
- |
  gluttonize
- |
  gluttonous
- |
  gluttonously
- |
  gluttony
- |
  glycerin
- |
  glycerine
- |
  glycerol
- |
  glycogen
- |
  glycogenic
- |
  Glyndwr
- |
  glyph
- |
  glyphic
- |
  glyptic
- |
  gnarl
- |
  gnarled
- |
  gnarly
- |
  gnash
- |
  gnathic
- |
  gnawer
- |
  gnawing
- |
  gneiss
- |
  gnocchi
- |
  gnome
- |
  gnomic
- |
  gnomically
- |
  gnomish
- |
  gnomon
- |
  gnomonic
- |
  gnosis
- |
  Gnostic
- |
  gnostic
- |
  Gnosticism
- |
  goalie
- |
  goalkeeper
- |
  goalkeeping
- |
  goalpost
- |
  goaltender
- |
  goatee
- |
  goatherd
- |
  goatish
- |
  goatskin
- |
  gobbet
- |
  gobble
- |
  gobbledegook
- |
  gobbledygook
- |
  gobbler
- |
  goblet
- |
  goblin
- |
  Godard
- |
  godchild
- |
  godchildren
- |
  goddammit
- |
  goddamn
- |
  goddamned
- |
  Goddard
- |
  goddaughter
- |
  goddess
- |
  godfather
- |
  godforsaken
- |
  Godfrey
- |
  Godhead
- |
  godhead
- |
  godhood
- |
  Godiva
- |
  godless
- |
  godlessly
- |
  godlessness
- |
  Godlike
- |
  godlike
- |
  godliness
- |
  godly
- |
  godmother
- |
  godparent
- |
  godsend
- |
  godson
- |
  Godspeed
- |
  Godthaab
- |
  Godthab
- |
  Godunov
- |
  Godwin
- |
  Goebbels
- |
  Goering
- |
  Goethals
- |
  Goethe
- |
  gofer
- |
  goggle
- |
  goggles
- |
  goggly
- |
  Gogol
- |
  Goiania
- |
  going
- |
  goiter
- |
  goitre
- |
  goitrous
- |
  Golconda
- |
  Goldberg
- |
  goldbrick
- |
  goldbricker
- |
  golden
- |
  goldenrod
- |
  goldfinch
- |
  goldfish
- |
  Goldilocks
- |
  Golding
- |
  Goldman
- |
  goldmine
- |
  Goldsmith
- |
  goldsmith
- |
  Goldwater
- |
  Goldwyn
- |
  golem
- |
  golfer
- |
  golfing
- |
  Golgotha
- |
  Goliath
- |
  golly
- |
  Gomel
- |
  Gomorrah
- |
  Gompers
- |
  gonad
- |
  gonadal
- |
  gonadic
- |
  gonadotropic
- |
  gonadotropin
- |
  gondola
- |
  gondolier
- |
  goner
- |
  gonfalon
- |
  gonfalonier
- |
  gonif
- |
  goniff
- |
  gonna
- |
  gonococcal
- |
  gonococci
- |
  gonococcus
- |
  gonorrhea
- |
  gonorrheal
- |
  gonorrhoea
- |
  gonzo
- |
  goober
- |
  goodby
- |
  goodbye
- |
  goodhearted
- |
  goodhumored
- |
  goodie
- |
  goodish
- |
  goodliness
- |
  goodly
- |
  Goodman
- |
  goodman
- |
  goodness
- |
  goodnight
- |
  goods
- |
  goodwife
- |
  goodwill
- |
  goody
- |
  Goodyear
- |
  gooey
- |
  goofball
- |
  goofily
- |
  goofiness
- |
  goofy
- |
  googol
- |
  goose
- |
  gooseberry
- |
  goosebumps
- |
  gooseflesh
- |
  gooseneck
- |
  goosenecked
- |
  Gopher
- |
  gopher
- |
  Gorbachev
- |
  Gordimer
- |
  Gordon
- |
  gored
- |
  Gorgas
- |
  gorge
- |
  gorgeous
- |
  gorgeously
- |
  gorgeousness
- |
  Gorgon
- |
  gorgon
- |
  Gorgonzola
- |
  gorilla
- |
  gorily
- |
  goriness
- |
  Gorki
- |
  Gorky
- |
  Gorlovka
- |
  gormandize
- |
  gormandizer
- |
  gormless
- |
  gormlessly
- |
  gormlessness
- |
  gorse
- |
  goshawk
- |
  gosling
- |
  Gospel
- |
  gospel
- |
  gossamer
- |
  gossamery
- |
  gossip
- |
  gossiper
- |
  gossipy
- |
  gotcha
- |
  Goteborg
- |
  Gothenburg
- |
  Gothic
- |
  gothic
- |
  Gothically
- |
  Gothicism
- |
  Gotland
- |
  gotta
- |
  gotten
- |
  gouache
- |
  Gouda
- |
  gouge
- |
  gouger
- |
  gouging
- |
  goulash
- |
  Gounod
- |
  gourami
- |
  gourd
- |
  gourde
- |
  gourmand
- |
  gourmandise
- |
  gourmandism
- |
  gourmet
- |
  goutiness
- |
  gouty
- |
  govern
- |
  governable
- |
  governance
- |
  governess
- |
  governing
- |
  Government
- |
  government
- |
  governmental
- |
  Governor
- |
  governor
- |
  governorship
- |
  goyim
- |
  goyish
- |
  grabber
- |
  grabby
- |
  Gracchus
- |
  Grace
- |
  grace
- |
  graceful
- |
  gracefully
- |
  gracefulness
- |
  graceless
- |
  gracelessly
- |
  Graces
- |
  graces
- |
  gracious
- |
  graciously
- |
  graciousness
- |
  grackle
- |
  gradate
- |
  gradation
- |
  gradational
- |
  grade
- |
  grader
- |
  gradient
- |
  gradual
- |
  gradualism
- |
  gradually
- |
  graduate
- |
  graduated
- |
  graduation
- |
  graduator
- |
  graffiti
- |
  graffitist
- |
  graffito
- |
  graft
- |
  grafter
- |
  Graham
- |
  graham
- |
  Grahame
- |
  Grail
- |
  grail
- |
  grain
- |
  grained
- |
  graininess
- |
  grainy
- |
  grammar
- |
  grammarian
- |
  grammatical
- |
  gramme
- |
  Grammy
- |
  gramophone
- |
  Grampian
- |
  grampus
- |
  Granada
- |
  granary
- |
  grand
- |
  grandam
- |
  grandame
- |
  grandchild
- |
  granddad
- |
  grandee
- |
  grandeur
- |
  grandfather
- |
  grandiose
- |
  grandiosely
- |
  grandiosity
- |
  grandly
- |
  grandma
- |
  grandmaster
- |
  grandmother
- |
  grandness
- |
  grandpa
- |
  grandparent
- |
  grandson
- |
  grandstand
- |
  grandstander
- |
  Grange
- |
  grange
- |
  granger
- |
  granite
- |
  graniteware
- |
  granitic
- |
  granitoid
- |
  grannie
- |
  granny
- |
  granola
- |
  Grant
- |
  grant
- |
  grantee
- |
  granter
- |
  grantor
- |
  granular
- |
  granularity
- |
  granulate
- |
  granulated
- |
  granulation
- |
  granulative
- |
  granule
- |
  Granville
- |
  grape
- |
  grapefruit
- |
  grapeshot
- |
  grapevine
- |
  graph
- |
  graphic
- |
  graphical
- |
  graphically
- |
  graphicness
- |
  graphics
- |
  graphite
- |
  graphitic
- |
  graphologist
- |
  graphology
- |
  grapnel
- |
  grapple
- |
  grappler
- |
  grasp
- |
  graspable
- |
  grasping
- |
  graspingly
- |
  Grass
- |
  grass
- |
  grasshopper
- |
  grassland
- |
  grassroots
- |
  grassy
- |
  grate
- |
  grated
- |
  grateful
- |
  gratefully
- |
  gratefulness
- |
  grater
- |
  Gratian
- |
  gratified
- |
  gratifier
- |
  gratify
- |
  gratifying
- |
  gratifyingly
- |
  grating
- |
  gratingly
- |
  gratis
- |
  gratitude
- |
  gratuitous
- |
  gratuitously
- |
  gratuity
- |
  gravamen
- |
  gravamina
- |
  grave
- |
  gravel
- |
  graveled
- |
  gravelly
- |
  gravely
- |
  graven
- |
  graveness
- |
  graver
- |
  Graves
- |
  graveside
- |
  gravestone
- |
  graveyard
- |
  gravid
- |
  gravidity
- |
  gravimeter
- |
  gravimetric
- |
  gravitas
- |
  gravitate
- |
  gravitater
- |
  gravitation
- |
  gravitative
- |
  graviton
- |
  gravity
- |
  gravure
- |
  gravy
- |
  graybeard
- |
  grayish
- |
  grayling
- |
  grayness
- |
  graze
- |
  grazed
- |
  grazer
- |
  grease
- |
  greaseless
- |
  greasepaint
- |
  greasewood
- |
  greasily
- |
  greasiness
- |
  greasy
- |
  great
- |
  greatcoat
- |
  greater
- |
  greathearted
- |
  greatly
- |
  greatness
- |
  grebe
- |
  Grecian
- |
  Greco
- |
  Greece
- |
  greed
- |
  greedily
- |
  greediness
- |
  greedy
- |
  Greek
- |
  Greeley
- |
  Green
- |
  green
- |
  greenback
- |
  greenbelt
- |
  Greene
- |
  greenery
- |
  greengrocer
- |
  greenhorn
- |
  greenhouse
- |
  greenish
- |
  Greenland
- |
  Greenlander
- |
  Greenlandic
- |
  greenly
- |
  greenmail
- |
  greenmailer
- |
  greenness
- |
  Greenpeace
- |
  greenroom
- |
  greens
- |
  Greensboro
- |
  greensward
- |
  Greenwich
- |
  greenwood
- |
  greeny
- |
  Greer
- |
  greet
- |
  greeter
- |
  greeting
- |
  greetings
- |
  gregarious
- |
  gregariously
- |
  Gregg
- |
  Gregory
- |
  gremlin
- |
  Grenada
- |
  grenade
- |
  Grenadian
- |
  grenadier
- |
  grenadine
- |
  Grenadines
- |
  Grenoble
- |
  Grenville
- |
  Gresham
- |
  Greta
- |
  Gretchen
- |
  Gretzky
- |
  greyhound
- |
  greyness
- |
  griddle
- |
  griddlecake
- |
  gridiron
- |
  gridlock
- |
  gridlocked
- |
  grief
- |
  Grieg
- |
  grievance
- |
  grieve
- |
  griever
- |
  grievous
- |
  grievously
- |
  grievousness
- |
  griffin
- |
  Griffith
- |
  griffon
- |
  grift
- |
  grifter
- |
  grill
- |
  grille
- |
  grilling
- |
  grillwork
- |
  grimace
- |
  grimacingly
- |
  grime
- |
  griminess
- |
  Grimke
- |
  grimly
- |
  Grimm
- |
  grimness
- |
  grimy
- |
  Grinch
- |
  grind
- |
  grinder
- |
  grinding
- |
  grindingly
- |
  grindstone
- |
  gringo
- |
  grinner
- |
  gripe
- |
  griper
- |
  gripes
- |
  griping
- |
  grippe
- |
  gripper
- |
  gripping
- |
  grippingly
- |
  grippy
- |
  grisaille
- |
  Griselda
- |
  grisliness
- |
  grisly
- |
  grist
- |
  gristle
- |
  gristly
- |
  gristmill
- |
  grits
- |
  gritter
- |
  grittily
- |
  grittiness
- |
  gritty
- |
  grizzled
- |
  grizzly
- |
  groan
- |
  groat
- |
  groats
- |
  grocer
- |
  groceries
- |
  grocery
- |
  Grodno
- |
  groggily
- |
  grogginess
- |
  groggy
- |
  groin
- |
  grommet
- |
  Gromyko
- |
  Groningen
- |
  groom
- |
  groomer
- |
  grooming
- |
  groomsman
- |
  groove
- |
  grooviness
- |
  groovy
- |
  grope
- |
  groper
- |
  groping
- |
  gropingly
- |
  Gropius
- |
  grosbeak
- |
  groschen
- |
  grosgrain
- |
  gross
- |
  grosses
- |
  grossly
- |
  grossness
- |
  Grosz
- |
  grosz
- |
  groszy
- |
  grotesque
- |
  grotesquely
- |
  grotesquery
- |
  grotto
- |
  grouch
- |
  grouchily
- |
  grouchiness
- |
  grouchy
- |
  ground
- |
  grounder
- |
  groundhog
- |
  grounding
- |
  groundless
- |
  groundlessly
- |
  groundling
- |
  grounds
- |
  groundswell
- |
  groundwater
- |
  groundwork
- |
  group
- |
  grouper
- |
  groupie
- |
  grouping
- |
  groupthink
- |
  groupware
- |
  grouse
- |
  grouser
- |
  grout
- |
  grouter
- |
  grove
- |
  grovel
- |
  groveler
- |
  grovelingly
- |
  groveller
- |
  Grover
- |
  grower
- |
  growl
- |
  growler
- |
  growly
- |
  grown
- |
  grownup
- |
  growth
- |
  Grozny
- |
  grubber
- |
  grubbily
- |
  grubbiness
- |
  grubby
- |
  grubstake
- |
  grudge
- |
  grudger
- |
  grudging
- |
  grudgingly
- |
  grudgingness
- |
  gruel
- |
  grueling
- |
  gruelingly
- |
  gruelling
- |
  gruesome
- |
  gruesomely
- |
  gruesomeness
- |
  gruff
- |
  gruffly
- |
  gruffness
- |
  grumble
- |
  grumbler
- |
  grumbly
- |
  grump
- |
  grumpily
- |
  grumpiness
- |
  grumps
- |
  grumpy
- |
  grunge
- |
  grunginess
- |
  grungy
- |
  grunion
- |
  grunt
- |
  grunter
- |
  Gruyere
- |
  gryphon
- |
  guacamole
- |
  Guadalajara
- |
  Guadalcanal
- |
  Guadalquivir
- |
  Guadalupe
- |
  Guadeloupe
- |
  Guallatiri
- |
  Guamanian
- |
  guanabana
- |
  Guanajuato
- |
  Guangzhou
- |
  guanine
- |
  guano
- |
  Guantanamo
- |
  Guarani
- |
  guarani
- |
  guarantee
- |
  guaranteed
- |
  guarantor
- |
  guaranty
- |
  guard
- |
  guarded
- |
  guardedly
- |
  guardedness
- |
  guarder
- |
  guardhouse
- |
  guardian
- |
  guardianship
- |
  guardrail
- |
  guardroom
- |
  guardsman
- |
  Guarneri
- |
  Guatemala
- |
  Guatemalan
- |
  guava
- |
  Guayaquil
- |
  Guenevere
- |
  guerdon
- |
  guerilla
- |
  Guernsey
- |
  Guerrero
- |
  guerrilla
- |
  guess
- |
  guesser
- |
  guesstimate
- |
  guesswork
- |
  guest
- |
  guesthouse
- |
  Guevara
- |
  guffaw
- |
  Guiana
- |
  Guianan
- |
  guidable
- |
  guidance
- |
  guide
- |
  guidebook
- |
  guideline
- |
  guidelines
- |
  guidepost
- |
  guider
- |
  guidon
- |
  guild
- |
  guilder
- |
  guildhall
- |
  guile
- |
  guileful
- |
  guilefully
- |
  guileless
- |
  guilelessly
- |
  guillotine
- |
  guilt
- |
  guiltily
- |
  guiltiness
- |
  guiltless
- |
  guiltlessly
- |
  guilty
- |
  Guinea
- |
  guinea
- |
  Guinean
- |
  Guinevere
- |
  Guinness
- |
  guise
- |
  guitar
- |
  guitarist
- |
  Guiyang
- |
  Guizot
- |
  Gujarati
- |
  Gujranwala
- |
  Gulag
- |
  gulag
- |
  gulch
- |
  gulden
- |
  gulfweed
- |
  Gullah
- |
  gullet
- |
  gullibility
- |
  gullible
- |
  gullibly
- |
  gully
- |
  gulper
- |
  Gumbo
- |
  gumbo
- |
  gumdrop
- |
  gummed
- |
  gumminess
- |
  gummy
- |
  gumption
- |
  gumshoe
- |
  gunboat
- |
  guncotton
- |
  gunfight
- |
  gunfighter
- |
  gunfire
- |
  gunky
- |
  gunlock
- |
  gunman
- |
  gunmetal
- |
  gunned
- |
  gunnel
- |
  gunner
- |
  gunnery
- |
  gunny
- |
  gunnysack
- |
  gunplay
- |
  gunpoint
- |
  gunpowder
- |
  gunrunner
- |
  gunrunning
- |
  gunsel
- |
  gunship
- |
  gunshot
- |
  gunslinger
- |
  gunsmith
- |
  gunwale
- |
  guppy
- |
  gurgle
- |
  gurgling
- |
  gurglingly
- |
  Gurkha
- |
  gurney
- |
  gusher
- |
  gushily
- |
  gushiness
- |
  gushing
- |
  gushy
- |
  gusset
- |
  gussie
- |
  gussy
- |
  gustatorily
- |
  gustatory
- |
  Gustavus
- |
  gustily
- |
  gustiness
- |
  gusto
- |
  gusty
- |
  Gutenberg
- |
  Guthrie
- |
  gutless
- |
  gutlessness
- |
  gutsily
- |
  gutsiness
- |
  gutsy
- |
  gutter
- |
  guttersnipe
- |
  guttural
- |
  gutturally
- |
  gutty
- |
  Guyana
- |
  Guyanese
- |
  guzzle
- |
  guzzler
- |
  Gwalior
- |
  Gwendoline
- |
  Gwendolyn
- |
  Gwent
- |
  Gwynedd
- |
  Gyandzha
- |
  gymkhana
- |
  gymnasia
- |
  gymnasial
- |
  gymnasium
- |
  gymnast
- |
  gymnastic
- |
  gymnastics
- |
  gymnosperm
- |
  gymnospermy
- |
  gynaecology
- |
  gynecologic
- |
  gynecologist
- |
  gynecology
- |
  gypper
- |
  gypster
- |
  gypsum
- |
  Gypsy
- |
  gypsy
- |
  gypsyish
- |
  gyrate
- |
  gyration
- |
  gyrator
- |
  gyratory
- |
  gyrfalcon
- |
  gyrocompass
- |
  gyros
- |
  gyroscope
- |
  gyroscopic
- |
  Haarlem
- |
  Habacuc
- |
  Habakkuk
- |
  habanera
- |
  haberdasher
- |
  haberdashery
- |
  habiliment
- |
  habiliments
- |
  habilitate
- |
  habilitation
- |
  habit
- |
  habitability
- |
  habitable
- |
  habitably
- |
  habitant
- |
  habitat
- |
  habitation
- |
  habitual
- |
  habitually
- |
  habitualness
- |
  habituate
- |
  habituation
- |
  habitude
- |
  habitue
- |
  Habsburg
- |
  hacek
- |
  hacienda
- |
  hackamore
- |
  hacker
- |
  hackery
- |
  hackie
- |
  hacking
- |
  hackle
- |
  hackles
- |
  hackman
- |
  Hackney
- |
  hackney
- |
  hackneyed
- |
  hacksaw
- |
  hackwork
- |
  haddock
- |
  Hadean
- |
  Hades
- |
  hades
- |
  hadji
- |
  Hadrian
- |
  hadron
- |
  hadrosaur
- |
  hadst
- |
  haecceity
- |
  haemoglobin
- |
  haemophiliac
- |
  haemorrhage
- |
  haemorrhoid
- |
  hafnium
- |
  Hagar
- |
  Haggai
- |
  haggard
- |
  haggardly
- |
  haggardness
- |
  haggis
- |
  haggish
- |
  haggle
- |
  haggler
- |
  haggling
- |
  Hagiographa
- |
  hagiographer
- |
  hagiographic
- |
  hagiography
- |
  Hague
- |
  hahnium
- |
  Haida
- |
  Haidarabad
- |
  Haifa
- |
  Haikou
- |
  haiku
- |
  hailer
- |
  hailstone
- |
  hailstorm
- |
  Haiphong
- |
  hairball
- |
  hairbreadth
- |
  hairbrush
- |
  haircloth
- |
  haircut
- |
  haircutter
- |
  haircutting
- |
  hairdo
- |
  hairdresser
- |
  hairdressing
- |
  hairdryer
- |
  haired
- |
  hairiness
- |
  hairless
- |
  hairlike
- |
  hairline
- |
  hairnet
- |
  hairpiece
- |
  hairpin
- |
  hairsbreadth
- |
  hairsplitter
- |
  hairspring
- |
  hairstyle
- |
  hairstyling
- |
  hairstylist
- |
  hairweaving
- |
  hairy
- |
  Haiti
- |
  Haitian
- |
  hajji
- |
  Hakluyt
- |
  halal
- |
  halala
- |
  halberd
- |
  halbert
- |
  halcyon
- |
  haleness
- |
  haler
- |
  Haley
- |
  halfback
- |
  halfcocked
- |
  halfhearted
- |
  halfpence
- |
  halfpenny
- |
  halftime
- |
  halftone
- |
  halftrack
- |
  halfway
- |
  halfwit
- |
  halfwitted
- |
  halibut
- |
  halide
- |
  Halifax
- |
  halite
- |
  halitosis
- |
  Halle
- |
  halleluiah
- |
  hallelujah
- |
  Halley
- |
  halliard
- |
  hallmark
- |
  hallmarked
- |
  hallo
- |
  halloo
- |
  hallow
- |
  hallowed
- |
  Halloween
- |
  hallower
- |
  hallucinant
- |
  hallucinate
- |
  hallucinator
- |
  hallucinogen
- |
  hallway
- |
  halocarbon
- |
  halogen
- |
  halogenous
- |
  Halsey
- |
  Halsingborg
- |
  halter
- |
  halting
- |
  haltingly
- |
  halvah
- |
  halve
- |
  halvers
- |
  halves
- |
  halyard
- |
  Hamadan
- |
  Hamadryad
- |
  hamadryad
- |
  hamadryades
- |
  Hamah
- |
  Hamal
- |
  Hamamatsu
- |
  hamartia
- |
  Hamas
- |
  Hamburg
- |
  hamburg
- |
  Hamburger
- |
  hamburger
- |
  Hamhung
- |
  Hamilton
- |
  Hamiltonian
- |
  Hamite
- |
  Hamitic
- |
  Hamlet
- |
  hamlet
- |
  Hammarskjold
- |
  Hammer
- |
  hammer
- |
  hammerer
- |
  hammerhead
- |
  hammering
- |
  hammerlock
- |
  Hammersmith
- |
  Hammerstein
- |
  hammertoe
- |
  Hammett
- |
  hammock
- |
  Hammurabi
- |
  Hammurapi
- |
  hammy
- |
  hamper
- |
  hamperer
- |
  Hampshire
- |
  Hampton
- |
  hamster
- |
  hamstring
- |
  hamstrings
- |
  hamstrung
- |
  Hamsun
- |
  Hancock
- |
  handbag
- |
  handball
- |
  handbarrow
- |
  handbill
- |
  handbook
- |
  handbreadth
- |
  handcar
- |
  handcart
- |
  handclasp
- |
  handcraft
- |
  handcuff
- |
  handcuffs
- |
  handed
- |
  Handel
- |
  handful
- |
  handgun
- |
  handheld
- |
  handicap
- |
  handicapped
- |
  handicapper
- |
  handicraft
- |
  handicrafter
- |
  handily
- |
  handiness
- |
  handiwork
- |
  handkerchief
- |
  handle
- |
  handlebar
- |
  handlebars
- |
  handled
- |
  handler
- |
  handless
- |
  handling
- |
  handmade
- |
  handmaid
- |
  handmaiden
- |
  handoff
- |
  handout
- |
  handover
- |
  handpick
- |
  handpicked
- |
  handrail
- |
  hands
- |
  handsaw
- |
  handsel
- |
  handset
- |
  handsful
- |
  handshake
- |
  handsome
- |
  handsomely
- |
  handsomeness
- |
  handspring
- |
  handstand
- |
  handwork
- |
  handwoven
- |
  handwriting
- |
  handwritten
- |
  Handy
- |
  handy
- |
  handyman
- |
  hangar
- |
  Hangchou
- |
  Hangchow
- |
  hangdog
- |
  hanger
- |
  hanging
- |
  hangman
- |
  hangnail
- |
  hangout
- |
  hangover
- |
  hangup
- |
  Hangzhou
- |
  hanker
- |
  hankerer
- |
  hankering
- |
  hankie
- |
  hanky
- |
  Hanna
- |
  Hannah
- |
  Hannibal
- |
  Hannover
- |
  Hanoi
- |
  Hanover
- |
  Hansberry
- |
  hansel
- |
  hansom
- |
  Hanuka
- |
  Hanukah
- |
  Hanukkah
- |
  haole
- |
  haphazard
- |
  haphazardly
- |
  hapless
- |
  haplessly
- |
  haplessness
- |
  haploid
- |
  haply
- |
  happen
- |
  happening
- |
  happenstance
- |
  happily
- |
  happiness
- |
  happy
- |
  Hapsburg
- |
  harangue
- |
  haranguer
- |
  Harare
- |
  harass
- |
  harassed
- |
  harasser
- |
  harassingly
- |
  harassment
- |
  Harbin
- |
  harbinger
- |
  harbor
- |
  harborage
- |
  harborer
- |
  harbour
- |
  hardback
- |
  hardball
- |
  hardboard
- |
  hardbound
- |
  hardcore
- |
  hardcover
- |
  harden
- |
  hardener
- |
  hardening
- |
  hardhack
- |
  hardhat
- |
  hardheaded
- |
  hardheadedly
- |
  hardhearted
- |
  hardihood
- |
  hardily
- |
  hardiness
- |
  Harding
- |
  hardline
- |
  hardliner
- |
  hardly
- |
  hardness
- |
  hardpan
- |
  hardscrabble
- |
  hardship
- |
  hardstand
- |
  hardtack
- |
  hardtop
- |
  hardware
- |
  hardwired
- |
  hardwood
- |
  hardworking
- |
  Hardy
- |
  hardy
- |
  harebell
- |
  harebrained
- |
  harelip
- |
  harelipped
- |
  harem
- |
  Haringey
- |
  harken
- |
  Harlan
- |
  Harland
- |
  Harlem
- |
  Harlemite
- |
  Harlequin
- |
  harlequin
- |
  Harley
- |
  harlot
- |
  harlotry
- |
  Harlow
- |
  harmful
- |
  harmfully
- |
  harmfulness
- |
  harmless
- |
  harmlessly
- |
  harmlessness
- |
  Harmon
- |
  harmonic
- |
  harmonica
- |
  harmonically
- |
  harmonics
- |
  harmonious
- |
  harmoniously
- |
  harmonise
- |
  harmonium
- |
  harmonize
- |
  harmonizer
- |
  harmony
- |
  Harmsworth
- |
  harness
- |
  harnesser
- |
  Harold
- |
  harper
- |
  harpist
- |
  harpoon
- |
  harpooner
- |
  harpsichord
- |
  Harpy
- |
  harpy
- |
  harquebus
- |
  harridan
- |
  harried
- |
  harrier
- |
  Harriet
- |
  Harriett
- |
  Harriette
- |
  Harris
- |
  Harrisburg
- |
  Harrison
- |
  Harrow
- |
  harrow
- |
  harrowing
- |
  Harry
- |
  harry
- |
  harsh
- |
  harshen
- |
  harshly
- |
  harshness
- |
  Harte
- |
  hartebeest
- |
  Hartford
- |
  harvest
- |
  harvester
- |
  harvesting
- |
  Harvey
- |
  hashish
- |
  Hasid
- |
  Hasidic
- |
  Hasidim
- |
  Hasidism
- |
  Hassid
- |
  Hassidim
- |
  hassium
- |
  hassle
- |
  hassock
- |
  haste
- |
  hasten
- |
  hastily
- |
  hastiness
- |
  Hastings
- |
  hasty
- |
  hatbox
- |
  hatch
- |
  hatchback
- |
  hatcheck
- |
  hatcher
- |
  hatchery
- |
  hatchet
- |
  hatching
- |
  hatchling
- |
  hatchway
- |
  hated
- |
  hateful
- |
  hatefully
- |
  hatefulness
- |
  hater
- |
  Hathaway
- |
  hatred
- |
  Hatshepset
- |
  Hatshepsut
- |
  hatter
- |
  Hattie
- |
  hauberk
- |
  haughtily
- |
  haughtiness
- |
  haughty
- |
  haulage
- |
  hauler
- |
  haunch
- |
  haunches
- |
  haunt
- |
  haunted
- |
  haunter
- |
  haunting
- |
  hauntingly
- |
  Hauptmann
- |
  Hausa
- |
  hauteur
- |
  Havana
- |
  Havanan
- |
  Havarti
- |
  Havel
- |
  haven
- |
  Havering
- |
  haversack
- |
  haves
- |
  havoc
- |
  Hawaii
- |
  Hawaiian
- |
  Hawke
- |
  hawker
- |
  Hawking
- |
  hawkish
- |
  hawkishly
- |
  hawkishness
- |
  Hawks
- |
  hawkweed
- |
  hawser
- |
  hawthorn
- |
  Hawthorne
- |
  haycock
- |
  Haydn
- |
  Hayes
- |
  hayfork
- |
  hayloft
- |
  haymow
- |
  hayrick
- |
  hayseed
- |
  haystack
- |
  Hayward
- |
  haywire
- |
  hazard
- |
  hazardous
- |
  hazardously
- |
  Hazel
- |
  hazel
- |
  hazelnut
- |
  hazer
- |
  hazily
- |
  haziness
- |
  hazing
- |
  Hazlitt
- |
  headache
- |
  headachy
- |
  headband
- |
  headboard
- |
  headdress
- |
  headed
- |
  header
- |
  headfirst
- |
  headgear
- |
  headhunter
- |
  headhunting
- |
  headily
- |
  headiness
- |
  heading
- |
  headlamp
- |
  headland
- |
  headless
- |
  headlight
- |
  headline
- |
  headliner
- |
  headlock
- |
  headlong
- |
  headman
- |
  headmaster
- |
  headmistress
- |
  headphone
- |
  headphones
- |
  headpiece
- |
  headpin
- |
  headquarters
- |
  headrest
- |
  headroom
- |
  heads
- |
  headset
- |
  headship
- |
  headshrink
- |
  headshrinker
- |
  headsman
- |
  headstall
- |
  headstand
- |
  headstone
- |
  headstrong
- |
  headteacher
- |
  headwaiter
- |
  headwater
- |
  headwaters
- |
  headway
- |
  headwind
- |
  headword
- |
  headwork
- |
  headworker
- |
  heady
- |
  healable
- |
  healer
- |
  health
- |
  healthful
- |
  healthfully
- |
  healthily
- |
  healthiness
- |
  healthy
- |
  Heaney
- |
  heaped
- |
  heaping
- |
  heaps
- |
  heard
- |
  hearer
- |
  hearing
- |
  hearken
- |
  hearsay
- |
  hearse
- |
  Hearst
- |
  heart
- |
  heartache
- |
  heartbeat
- |
  heartbreak
- |
  heartbreaker
- |
  heartbroken
- |
  heartburn
- |
  hearted
- |
  hearten
- |
  heartened
- |
  heartening
- |
  heartfelt
- |
  hearth
- |
  hearthstone
- |
  heartily
- |
  heartiness
- |
  heartland
- |
  heartless
- |
  heartlessly
- |
  heartrending
- |
  heartsick
- |
  heartstrings
- |
  heartthrob
- |
  heartwarming
- |
  heartwood
- |
  hearty
- |
  heated
- |
  heatedly
- |
  heater
- |
  Heath
- |
  heath
- |
  heathen
- |
  heathendom
- |
  heathenish
- |
  heathenism
- |
  heathenry
- |
  Heather
- |
  heather
- |
  heathery
- |
  heathy
- |
  heating
- |
  heatproof
- |
  heatstroke
- |
  heave
- |
  Heaven
- |
  heaven
- |
  heavenliness
- |
  heavenly
- |
  heavens
- |
  heavenward
- |
  heavenwards
- |
  heaver
- |
  heaves
- |
  heavily
- |
  heaviness
- |
  heavy
- |
  heavyhearted
- |
  heavyish
- |
  heavyset
- |
  heavyweight
- |
  hebdomadal
- |
  hebetude
- |
  Hebraic
- |
  Hebraism
- |
  Hebraist
- |
  Hebraistic
- |
  Hebraistical
- |
  Hebrew
- |
  Hebrews
- |
  Hebridean
- |
  Hebrides
- |
  hecatomb
- |
  heckle
- |
  heckler
- |
  heckling
- |
  hectarage
- |
  hectare
- |
  hectic
- |
  hectically
- |
  hectogram
- |
  hectoliter
- |
  hectometer
- |
  Hector
- |
  hector
- |
  hectoring
- |
  hectoringly
- |
  Hecuba
- |
  hedge
- |
  hedgehog
- |
  hedgehop
- |
  hedger
- |
  hedgerow
- |
  hedonism
- |
  hedonist
- |
  hedonistic
- |
  heedful
- |
  heedfully
- |
  heedfulness
- |
  heedless
- |
  heedlessly
- |
  heedlessness
- |
  heehaw
- |
  heeled
- |
  heels
- |
  heftily
- |
  heftiness
- |
  hefty
- |
  Hegel
- |
  hegemonic
- |
  hegemonism
- |
  hegemonist
- |
  hegemony
- |
  Hegira
- |
  hegira
- |
  Heidegger
- |
  Heidelberg
- |
  Heidi
- |
  heifer
- |
  Heifetz
- |
  height
- |
  heighten
- |
  heights
- |
  Heilongjiang
- |
  Heilungkiang
- |
  Heine
- |
  heinous
- |
  heinously
- |
  heinousness
- |
  Heinz
- |
  heiress
- |
  heirloom
- |
  heirship
- |
  Heisenberg
- |
  heist
- |
  Hejira
- |
  Helaine
- |
  Helen
- |
  Helena
- |
  Helene
- |
  Helga
- |
  helical
- |
  helically
- |
  helices
- |
  helicopter
- |
  heliocentric
- |
  Heliopolis
- |
  Helios
- |
  heliotrope
- |
  heliport
- |
  helium
- |
  helix
- |
  hellbent
- |
  hellcat
- |
  hellebore
- |
  Hellene
- |
  Hellenic
- |
  Hellenism
- |
  Hellenist
- |
  Hellenistic
- |
  Hellenize
- |
  Hellenizer
- |
  Heller
- |
  Hellespont
- |
  hellgrammite
- |
  hellhole
- |
  hellion
- |
  hellish
- |
  hellishly
- |
  hellishness
- |
  Hellman
- |
  hello
- |
  helmet
- |
  helminth
- |
  helmsman
- |
  Helmut
- |
  Heloise
- |
  helot
- |
  helotage
- |
  helotism
- |
  helotry
- |
  helper
- |
  helpful
- |
  helpfully
- |
  helpfulness
- |
  helping
- |
  helpless
- |
  helplessly
- |
  helplessness
- |
  helpline
- |
  helpmate
- |
  helpmeet
- |
  Helsinki
- |
  helve
- |
  Helvetia
- |
  Helvetian
- |
  hematite
- |
  hematologic
- |
  hematologist
- |
  hematology
- |
  hematoma
- |
  hematomata
- |
  Hemings
- |
  Hemingway
- |
  hemisphere
- |
  hemispheric
- |
  hemline
- |
  hemlock
- |
  hemmer
- |
  hemodialyses
- |
  hemodialysis
- |
  hemoglobin
- |
  hemophilia
- |
  hemophiliac
- |
  hemorrhage
- |
  hemorrhagic
- |
  hemorrhaging
- |
  hemorrhoid
- |
  hemorrhoidal
- |
  hemorrhoids
- |
  hemostat
- |
  hemostatic
- |
  hempen
- |
  hemstitch
- |
  hence
- |
  henceforth
- |
  henceforward
- |
  henchman
- |
  hendiadys
- |
  Hendrix
- |
  henna
- |
  henotheism
- |
  henpeck
- |
  henpecked
- |
  Henrietta
- |
  Henry
- |
  henry
- |
  Henson
- |
  heparin
- |
  hepatic
- |
  hepatica
- |
  hepatitis
- |
  Hepburn
- |
  Hephaestus
- |
  heptagon
- |
  heptagonal
- |
  heptameter
- |
  heptathlon
- |
  Heracles
- |
  Heraclitean
- |
  Heraclitus
- |
  Heraklion
- |
  herald
- |
  heraldic
- |
  heraldically
- |
  heraldist
- |
  heraldry
- |
  Herat
- |
  herbaceous
- |
  herbage
- |
  herbal
- |
  herbalism
- |
  herbalist
- |
  herbaria
- |
  herbarium
- |
  Herbert
- |
  herbicidal
- |
  herbicide
- |
  herbivore
- |
  herbivorous
- |
  herby
- |
  Herculaneum
- |
  Herculean
- |
  herculean
- |
  Hercules
- |
  Herder
- |
  herder
- |
  herdsman
- |
  hereabout
- |
  hereabouts
- |
  hereafter
- |
  hereby
- |
  hereditarily
- |
  hereditary
- |
  heredity
- |
  Hereford
- |
  herein
- |
  hereof
- |
  hereon
- |
  heresy
- |
  heretic
- |
  heretical
- |
  heretically
- |
  hereto
- |
  heretofore
- |
  hereunder
- |
  hereunto
- |
  hereupon
- |
  herewith
- |
  heritability
- |
  heritable
- |
  heritably
- |
  heritage
- |
  Herman
- |
  Hermann
- |
  hermeneutic
- |
  Hermes
- |
  Hermetic
- |
  hermetic
- |
  hermetical
- |
  hermetically
- |
  hermeticism
- |
  Hermine
- |
  hermit
- |
  Hermitage
- |
  hermitage
- |
  hermitic
- |
  Hermosillo
- |
  hernia
- |
  herniae
- |
  hernial
- |
  herniate
- |
  herniation
- |
  Herod
- |
  Herodotus
- |
  heroic
- |
  heroical
- |
  heroically
- |
  heroics
- |
  heroin
- |
  heroine
- |
  heroism
- |
  heron
- |
  herpes
- |
  herpetic
- |
  herpetologic
- |
  herpetology
- |
  Herren
- |
  Herrick
- |
  herring
- |
  herringbone
- |
  Herschel
- |
  herself
- |
  Hershel
- |
  Hertford
- |
  hertz
- |
  Herzegovina
- |
  Herzl
- |
  Heshvan
- |
  Heshwan
- |
  Hesiod
- |
  hesitance
- |
  hesitancy
- |
  hesitant
- |
  hesitantly
- |
  hesitate
- |
  hesitatingly
- |
  hesitation
- |
  Hesse
- |
  Hester
- |
  Hestia
- |
  heteroclite
- |
  heteroclitic
- |
  heterodox
- |
  heterodoxy
- |
  heterogenous
- |
  heteronym
- |
  heteronymic
- |
  heteronymous
- |
  heterosexual
- |
  heterotroph
- |
  heterotrophy
- |
  heuristic
- |
  heuristics
- |
  hewer
- |
  hexadecimal
- |
  hexagon
- |
  hexagonal
- |
  hexagonally
- |
  hexagram
- |
  hexameter
- |
  hexametric
- |
  hexametrical
- |
  hexer
- |
  heyday
- |
  Heyerdahl
- |
  Hezbollah
- |
  Hialeah
- |
  hiatal
- |
  hiatus
- |
  Hiawatha
- |
  hibachi
- |
  hibernate
- |
  hibernation
- |
  hibernator
- |
  Hibernia
- |
  Hibernian
- |
  hibiscus
- |
  hiccough
- |
  hiccoughs
- |
  hiccup
- |
  hiccups
- |
  hickey
- |
  Hickok
- |
  hickory
- |
  Hidalgo
- |
  hidalgo
- |
  hidden
- |
  hideaway
- |
  hidebound
- |
  hideous
- |
  hideously
- |
  hideousness
- |
  hideout
- |
  hider
- |
  hiding
- |
  hidrosis
- |
  hidrotic
- |
  hierarchal
- |
  hierarchic
- |
  hierarchical
- |
  hierarchize
- |
  hierarchy
- |
  hieratic
- |
  hieratically
- |
  hierocracy
- |
  hierocratic
- |
  hieroglyph
- |
  hieroglyphic
- |
  hierophant
- |
  hifalutin
- |
  Higashiosaka
- |
  highball
- |
  highborn
- |
  highboy
- |
  highbred
- |
  highbrow
- |
  highbrowed
- |
  highbrowism
- |
  highchair
- |
  highfalutin
- |
  highfaluting
- |
  highhanded
- |
  highhandedly
- |
  highjack
- |
  Highland
- |
  highland
- |
  Highlander
- |
  highlander
- |
  Highlands
- |
  highlands
- |
  highlight
- |
  highlighter
- |
  highly
- |
  Highness
- |
  highness
- |
  highroad
- |
  hightail
- |
  hightest
- |
  highway
- |
  highwayman
- |
  hijack
- |
  hijacker
- |
  hijacking
- |
  hijinks
- |
  Hijra
- |
  hiker
- |
  hiking
- |
  hilarious
- |
  hilariously
- |
  hilarity
- |
  Hilary
- |
  Hilda
- |
  Hildegard
- |
  Hildegarde
- |
  Hillary
- |
  hillbilly
- |
  hilliness
- |
  Hillingdon
- |
  hillock
- |
  hillside
- |
  hilltop
- |
  hilly
- |
  Hilton
- |
  Hilwan
- |
  Himalaya
- |
  Himalayan
- |
  Himalayas
- |
  Himmler
- |
  himself
- |
  Hindemith
- |
  Hindenburg
- |
  hinder
- |
  hinderer
- |
  hindermost
- |
  Hindi
- |
  hindmost
- |
  hindquarter
- |
  hindquarters
- |
  hindrance
- |
  hindsight
- |
  Hindu
- |
  Hinduism
- |
  Hindustan
- |
  Hindustani
- |
  Hines
- |
  hinge
- |
  hinged
- |
  hinter
- |
  hinterland
- |
  hinterlands
- |
  hipbone
- |
  hiphop
- |
  hipness
- |
  hipped
- |
  hippie
- |
  hippiedom
- |
  hippo
- |
  hippocampi
- |
  hippocampus
- |
  Hippocrates
- |
  Hippocratic
- |
  hippodrome
- |
  hippopotami
- |
  hippopotamus
- |
  hippy
- |
  hipster
- |
  hiragana
- |
  Hiram
- |
  hircine
- |
  hireling
- |
  hirer
- |
  Hirohito
- |
  Hiroshima
- |
  hirsute
- |
  hirsuteness
- |
  Hispanic
- |
  Hispanicize
- |
  Hispaniola
- |
  hissing
- |
  histamine
- |
  histaminic
- |
  histogram
- |
  histologic
- |
  histological
- |
  histologist
- |
  histology
- |
  historian
- |
  historic
- |
  historical
- |
  historically
- |
  historicism
- |
  historicist
- |
  historicity
- |
  history
- |
  histrionic
- |
  histrionical
- |
  histrionics
- |
  hitch
- |
  Hitchcock
- |
  hitcher
- |
  hitchhike
- |
  hitchhiker
- |
  hitchhiking
- |
  hither
- |
  hitherto
- |
  Hitler
- |
  Hitlerian
- |
  hitter
- |
  Hittite
- |
  hives
- |
  Hmong
- |
  hoagie
- |
  hoagy
- |
  hoard
- |
  hoarded
- |
  hoarder
- |
  hoarding
- |
  hoarfrost
- |
  hoarily
- |
  hoariness
- |
  hoarse
- |
  hoarsely
- |
  hoarseness
- |
  hoary
- |
  hoaxer
- |
  Hobart
- |
  Hobbes
- |
  Hobbesian
- |
  hobble
- |
  hobbledehoy
- |
  hobbler
- |
  hobby
- |
  hobbyhorse
- |
  hobbyist
- |
  hobgoblin
- |
  hobnail
- |
  hobnailed
- |
  hobnob
- |
  hockey
- |
  Hockney
- |
  hockshop
- |
  hodgepodge
- |
  Hodgkin
- |
  hoecake
- |
  hoedown
- |
  Hoffa
- |
  hogan
- |
  Hogarth
- |
  Hogarthian
- |
  hogback
- |
  hogger
- |
  hoggish
- |
  hoggishly
- |
  hogshead
- |
  hogtie
- |
  hogwash
- |
  Hohhot
- |
  hoist
- |
  hoister
- |
  Hokan
- |
  hokey
- |
  Hokkaido
- |
  hokku
- |
  hokum
- |
  Holarctic
- |
  Holbein
- |
  holder
- |
  holding
- |
  holdings
- |
  holdout
- |
  holdover
- |
  holdup
- |
  holey
- |
  Holguin
- |
  Holiday
- |
  holiday
- |
  holidaymaker
- |
  holidays
- |
  holily
- |
  Holiness
- |
  holiness
- |
  Holinshed
- |
  holism
- |
  holist
- |
  holistic
- |
  holistically
- |
  Holland
- |
  Hollander
- |
  holler
- |
  Hollis
- |
  hollow
- |
  holloware
- |
  hollowly
- |
  hollowness
- |
  hollowware
- |
  Holly
- |
  holly
- |
  hollyhock
- |
  Hollywood
- |
  Holmes
- |
  holmium
- |
  Holocaust
- |
  holocaust
- |
  Holocene
- |
  hologram
- |
  holograph
- |
  holographic
- |
  holography
- |
  holophrase
- |
  holophrasis
- |
  holophrastic
- |
  Holst
- |
  Holstein
- |
  holster
- |
  holstered
- |
  holystone
- |
  homage
- |
  hombre
- |
  Homburg
- |
  homburg
- |
  homebody
- |
  homeboy
- |
  homebred
- |
  homecoming
- |
  homegirl
- |
  homegrown
- |
  homeland
- |
  homeless
- |
  homelessness
- |
  homelike
- |
  homeliness
- |
  homely
- |
  homemade
- |
  homemaker
- |
  homemaking
- |
  homeopath
- |
  homeopathic
- |
  homeopathist
- |
  homeopathy
- |
  homeostases
- |
  homeostasis
- |
  homeostatic
- |
  homeotherm
- |
  homeowner
- |
  homepage
- |
  Homer
- |
  homer
- |
  Homeric
- |
  homeroom
- |
  homeschool
- |
  homeschooler
- |
  homesick
- |
  homesickness
- |
  homespun
- |
  homestead
- |
  homesteader
- |
  homesteading
- |
  homestretch
- |
  hometown
- |
  homeward
- |
  homewards
- |
  homework
- |
  homey
- |
  homeyness
- |
  homicidal
- |
  Homicide
- |
  homicide
- |
  homiletic
- |
  homiletics
- |
  homilist
- |
  homily
- |
  hominess
- |
  hominid
- |
  hominoid
- |
  hominy
- |
  homoeopathy
- |
  homoerotic
- |
  homogeneity
- |
  homogeneous
- |
  homogenize
- |
  homogenized
- |
  homogenizer
- |
  homogenous
- |
  homogeny
- |
  homograph
- |
  homographic
- |
  homolog
- |
  homologous
- |
  homologue
- |
  homology
- |
  homonym
- |
  homonymic
- |
  homonymous
- |
  homonymy
- |
  homophobe
- |
  homophobia
- |
  homophobic
- |
  homophone
- |
  homophonic
- |
  homophonous
- |
  homophony
- |
  homosexual
- |
  honcho
- |
  Hondo
- |
  Honduran
- |
  Honduranean
- |
  Honduranian
- |
  Honduras
- |
  Honecker
- |
  honer
- |
  honest
- |
  honestly
- |
  honesty
- |
  honey
- |
  honeybee
- |
  honeycomb
- |
  honeycombed
- |
  honeydew
- |
  honeyed
- |
  honeylocust
- |
  honeymoon
- |
  honeymooner
- |
  honeysuckle
- |
  Honiara
- |
  honied
- |
  honker
- |
  honky
- |
  Honolulu
- |
  Honor
- |
  honor
- |
  Honorable
- |
  honorable
- |
  honorably
- |
  honoraria
- |
  honorarily
- |
  honorarium
- |
  honorary
- |
  honoree
- |
  honorer
- |
  honorific
- |
  honors
- |
  honour
- |
  honourable
- |
  honourably
- |
  honoured
- |
  Honshu
- |
  hooch
- |
  hooded
- |
  hoodlum
- |
  hoodlumism
- |
  hoodoo
- |
  hoodwink
- |
  hoodwinker
- |
  hooey
- |
  hoofed
- |
  Hooghly
- |
  hooka
- |
  hookah
- |
  Hooke
- |
  hooked
- |
  Hooker
- |
  hooker
- |
  hookey
- |
  hookup
- |
  hookworm
- |
  hooky
- |
  hooligan
- |
  hooliganism
- |
  hoopla
- |
  hoops
- |
  hooray
- |
  hoosegow
- |
  Hoosier
- |
  hootenanny
- |
  hooter
- |
  Hoover
- |
  hoover
- |
  hoovering
- |
  Hooverville
- |
  hooves
- |
  hopeful
- |
  hopefully
- |
  hopefulness
- |
  hopeless
- |
  hopelessly
- |
  hopelessness
- |
  hophead
- |
  Hopkins
- |
  Hopper
- |
  hopper
- |
  hopsack
- |
  hopsacking
- |
  hopscotch
- |
  Horace
- |
  horah
- |
  Horatian
- |
  Horatio
- |
  horde
- |
  horehound
- |
  horizon
- |
  horizons
- |
  horizontal
- |
  horizontally
- |
  Horlivka
- |
  hormonal
- |
  hormonally
- |
  hormone
- |
  Hormuz
- |
  hornblende
- |
  hornbook
- |
  Horne
- |
  horned
- |
  hornet
- |
  horniness
- |
  hornless
- |
  hornlike
- |
  hornpipe
- |
  horny
- |
  horologer
- |
  horologic
- |
  horological
- |
  horologist
- |
  Horologium
- |
  horology
- |
  horoscope
- |
  Horowitz
- |
  horrendous
- |
  horrendously
- |
  horrible
- |
  horribleness
- |
  horribly
- |
  horrid
- |
  horridly
- |
  horridness
- |
  horrific
- |
  horrifically
- |
  horrified
- |
  horrify
- |
  horrifying
- |
  horrifyingly
- |
  horror
- |
  horse
- |
  horseback
- |
  horseflesh
- |
  horsefly
- |
  horsehair
- |
  horsehide
- |
  horselaugh
- |
  horseless
- |
  horseman
- |
  horsemanship
- |
  horseplay
- |
  horseplayer
- |
  horsepower
- |
  horseracing
- |
  horseradish
- |
  horseshoe
- |
  horseshoer
- |
  horseshoes
- |
  horsetail
- |
  horsewhip
- |
  horsewoman
- |
  horsey
- |
  horsily
- |
  horsiness
- |
  horsy
- |
  hortation
- |
  hortative
- |
  hortatory
- |
  Hortense
- |
  horticulture
- |
  Horus
- |
  hosanna
- |
  hosannah
- |
  Hosea
- |
  hosiery
- |
  hospice
- |
  hospitable
- |
  hospitably
- |
  hospital
- |
  Hospitalet
- |
  hospitalise
- |
  hospitality
- |
  hospitalize
- |
  hosta
- |
  hostage
- |
  hostel
- |
  hosteler
- |
  hostelry
- |
  hostess
- |
  hostile
- |
  hostilely
- |
  hostilities
- |
  hostility
- |
  hostler
- |
  hotbed
- |
  hotblooded
- |
  hotbox
- |
  hotcake
- |
  hotchpotch
- |
  hotdog
- |
  hotel
- |
  hotelier
- |
  hotfoot
- |
  hothead
- |
  hotheaded
- |
  hotheadedly
- |
  hothouse
- |
  hotline
- |
  hotlink
- |
  hotly
- |
  hotness
- |
  hotplate
- |
  hotshot
- |
  hotspot
- |
  Hottentot
- |
  Houdini
- |
  hound
- |
  hounder
- |
  Hounslow
- |
  hourglass
- |
  houri
- |
  hourly
- |
  hours
- |
  House
- |
  house
- |
  houseboat
- |
  housebound
- |
  houseboy
- |
  housebreak
- |
  housebreaker
- |
  housebroke
- |
  housebroken
- |
  houseclean
- |
  housecoat
- |
  housefly
- |
  houseful
- |
  household
- |
  householder
- |
  househusband
- |
  housekeeper
- |
  housekeeping
- |
  houselights
- |
  housemaid
- |
  housemother
- |
  houseplant
- |
  housetop
- |
  housewares
- |
  housewarming
- |
  housewife
- |
  housewifely
- |
  housewifery
- |
  housewives
- |
  housework
- |
  houseworker
- |
  housing
- |
  Housman
- |
  Houston
- |
  Houstonian
- |
  hovel
- |
  hover
- |
  hovercraft
- |
  Howard
- |
  howbeit
- |
  howdah
- |
  howdy
- |
  Howell
- |
  Howells
- |
  however
- |
  howitzer
- |
  howler
- |
  howling
- |
  Howrah
- |
  howsoever
- |
  Hoxha
- |
  hoyden
- |
  hoydenish
- |
  Hoyle
- |
  hryvnia
- |
  Huang
- |
  huarache
- |
  huaraches
- |
  Huascaran
- |
  Hubble
- |
  hubbub
- |
  hubby
- |
  hubcap
- |
  Hubert
- |
  Hubli
- |
  hubris
- |
  hubristic
- |
  huckleberry
- |
  huckster
- |
  hucksterism
- |
  Huddersfield
- |
  huddle
- |
  huddler
- |
  Hudson
- |
  huffily
- |
  huffiness
- |
  huffy
- |
  hugely
- |
  hugeness
- |
  hugger
- |
  Hughes
- |
  Hugli
- |
  Huguenot
- |
  Huhehot
- |
  hulking
- |
  hulky
- |
  hullaballoo
- |
  hullabaloo
- |
  huller
- |
  hullo
- |
  human
- |
  humane
- |
  humanely
- |
  humaneness
- |
  humanhood
- |
  Humanism
- |
  humanism
- |
  humanist
- |
  humanistic
- |
  humanitarian
- |
  humanities
- |
  humanity
- |
  humanization
- |
  humanize
- |
  humanizer
- |
  humankind
- |
  humanly
- |
  humanness
- |
  humanoid
- |
  Humberside
- |
  humble
- |
  humbled
- |
  humbleness
- |
  humbler
- |
  humbling
- |
  humbly
- |
  Humboldt
- |
  humbug
- |
  humbugger
- |
  humbuggery
- |
  humdinger
- |
  humdrum
- |
  humectant
- |
  humeral
- |
  humeri
- |
  humerus
- |
  humid
- |
  humidifier
- |
  humidify
- |
  humidity
- |
  humidly
- |
  humidor
- |
  humiliate
- |
  humiliated
- |
  humiliating
- |
  humiliation
- |
  humility
- |
  hummable
- |
  hummer
- |
  humming
- |
  hummingbird
- |
  hummock
- |
  hummocky
- |
  hummus
- |
  humongous
- |
  humor
- |
  humoresque
- |
  humorist
- |
  humorless
- |
  humorlessly
- |
  humorous
- |
  humorously
- |
  humorousness
- |
  humour
- |
  humpback
- |
  humpbacked
- |
  humped
- |
  Humperdinck
- |
  Humphrey
- |
  Humphry
- |
  humungous
- |
  humus
- |
  Humvee
- |
  Hunan
- |
  hunch
- |
  hunchback
- |
  hunchbacked
- |
  hunched
- |
  hundred
- |
  hundredfold
- |
  hundreds
- |
  hundredth
- |
  Hungarian
- |
  Hungary
- |
  hunger
- |
  hungover
- |
  hungrily
- |
  hungriness
- |
  hungry
- |
  hunker
- |
  hunkers
- |
  hunky
- |
  hunter
- |
  hunting
- |
  Huntington
- |
  huntress
- |
  huntsman
- |
  Huntsville
- |
  hurdle
- |
  hurdler
- |
  hurler
- |
  Huron
- |
  hurrah
- |
  hurray
- |
  hurricane
- |
  hurried
- |
  hurriedly
- |
  hurriedness
- |
  hurry
- |
  Hurston
- |
  hurtful
- |
  hurtfully
- |
  hurtfulness
- |
  hurtle
- |
  Husain
- |
  husband
- |
  husbander
- |
  husbandman
- |
  husbandry
- |
  hushed
- |
  husker
- |
  huskily
- |
  huskiness
- |
  husky
- |
  hussar
- |
  Hussein
- |
  Husserl
- |
  hussy
- |
  hustings
- |
  hustle
- |
  hustler
- |
  Huston
- |
  hutch
- |
  Hutchinson
- |
  Hutton
- |
  hutzpa
- |
  hutzpah
- |
  Huxley
- |
  huzza
- |
  huzzah
- |
  Hwang
- |
  hyacinth
- |
  hyaena
- |
  hybrid
- |
  hybridism
- |
  hybridity
- |
  hybridize
- |
  hybridizer
- |
  Hyderabad
- |
  Hydra
- |
  hydra
- |
  hydrangea
- |
  hydrant
- |
  hydratable
- |
  hydrate
- |
  hydrated
- |
  hydration
- |
  hydrator
- |
  hydraulic
- |
  hydraulics
- |
  hydro
- |
  hydrocarbon
- |
  hydrocephaly
- |
  hydrodynamic
- |
  hydrofoil
- |
  hydrogen
- |
  hydrogenate
- |
  hydrogenous
- |
  hydrographer
- |
  hydrographic
- |
  hydrography
- |
  hydrologic
- |
  hydrological
- |
  hydrologist
- |
  hydrology
- |
  hydrolyses
- |
  hydrolysis
- |
  hydrolyte
- |
  hydrolytic
- |
  hydrolyze
- |
  hydrometer
- |
  hydrometric
- |
  hydrometry
- |
  hydropathic
- |
  hydropathist
- |
  hydropathy
- |
  hydrophobia
- |
  hydrophobic
- |
  hydrophone
- |
  hydroplane
- |
  hydroponic
- |
  hydroponics
- |
  hydropower
- |
  hydrosphere
- |
  hydrostatic
- |
  hydrostatics
- |
  hydrotherapy
- |
  hydrothermal
- |
  hydrous
- |
  hydroxide
- |
  Hydrus
- |
  hyena
- |
  hygiene
- |
  hygienic
- |
  hygienically
- |
  hygienist
- |
  hygrometer
- |
  hygrometric
- |
  hygrometry
- |
  hygroscopic
- |
  hying
- |
  Hymen
- |
  hymen
- |
  hymenal
- |
  hymeneal
- |
  hymnal
- |
  hymnbook
- |
  hyper
- |
  hyperacid
- |
  hyperacidity
- |
  hyperactive
- |
  hyperbaric
- |
  hyperbola
- |
  hyperbolae
- |
  hyperbole
- |
  hyperbolic
- |
  hyperbolical
- |
  hyperbolism
- |
  hyperlink
- |
  hypermedia
- |
  hyperopia
- |
  hyperopic
- |
  hypersonic
- |
  hyperspace
- |
  hyperspatial
- |
  hypertension
- |
  hypertensive
- |
  hypertext
- |
  hyperthermia
- |
  hyperthyroid
- |
  hypertrophic
- |
  hypertrophy
- |
  hyphen
- |
  hyphenate
- |
  hyphenated
- |
  hyphenation
- |
  hypnagogic
- |
  hypnogogic
- |
  hypnoses
- |
  hypnosis
- |
  hypnotherapy
- |
  hypnotic
- |
  hypnotically
- |
  hypnotism
- |
  hypnotist
- |
  hypnotizable
- |
  hypnotize
- |
  hypnotizer
- |
  hypocenter
- |
  hypochondria
- |
  hypocrisy
- |
  hypocrite
- |
  hypocritical
- |
  hypodermic
- |
  hypoglycemia
- |
  hypoglycemic
- |
  hypostases
- |
  hypostasis
- |
  hypotension
- |
  hypotenuse
- |
  hypothalami
- |
  hypothalamic
- |
  hypothalamus
- |
  hypothermia
- |
  hypothermic
- |
  hypotheses
- |
  hypothesis
- |
  hypothesize
- |
  hypothetic
- |
  hypothetical
- |
  hypothyroid
- |
  hyraces
- |
  hyrax
- |
  hyssop
- |
  hysterectomy
- |
  hysteria
- |
  hysteric
- |
  hysterical
- |
  hysterically
- |
  hysterics
- |
  Iacocca
- |
  iambi
- |
  iambic
- |
  iambus
- |
  Ibadan
- |
  Ibague
- |
  Iberia
- |
  Iberian
- |
  ibices
- |
  ibidem
- |
  Ibiza
- |
  Ibsen
- |
  ibuprofen
- |
  Icarus
- |
  iceberg
- |
  iceboat
- |
  iceboater
- |
  iceboating
- |
  icebound
- |
  icebox
- |
  icebreaker
- |
  icebreaking
- |
  icecap
- |
  icehouse
- |
  Iceland
- |
  Icelander
- |
  Icelandic
- |
  iceman
- |
  Ichabod
- |
  ichor
- |
  ichorous
- |
  ichthyologic
- |
  ichthyology
- |
  ichthyosaur
- |
  icicle
- |
  icily
- |
  iciness
- |
  icing
- |
  ickiness
- |
  iconic
- |
  iconically
- |
  iconicity
- |
  iconoclasm
- |
  iconoclast
- |
  iconoclastic
- |
  ictus
- |
  Idaho
- |
  Idahoan
- |
  ideal
- |
  idealise
- |
  idealism
- |
  idealist
- |
  idealistic
- |
  idealization
- |
  idealize
- |
  idealized
- |
  idealizer
- |
  ideally
- |
  idealogy
- |
  ideate
- |
  ideated
- |
  ideation
- |
  ideational
- |
  identical
- |
  identically
- |
  identifiable
- |
  identifiably
- |
  identifier
- |
  identify
- |
  identity
- |
  ideogram
- |
  ideograph
- |
  ideographic
- |
  ideography
- |
  ideological
- |
  ideologist
- |
  ideologue
- |
  ideology
- |
  idiocy
- |
  idiographic
- |
  idiom
- |
  idiomatic
- |
  idiopathic
- |
  idiopathy
- |
  idiosyncrasy
- |
  idiot
- |
  idiotic
- |
  idiotically
- |
  idiotropic
- |
  idleness
- |
  idler
- |
  idolater
- |
  idolator
- |
  idolatrous
- |
  idolatrously
- |
  idolatry
- |
  idolization
- |
  idolize
- |
  idolizer
- |
  idyll
- |
  idyllic
- |
  idyllically
- |
  idyllist
- |
  idyllize
- |
  iffiness
- |
  igloo
- |
  Ignatius
- |
  igneous
- |
  ignitable
- |
  ignite
- |
  ignitible
- |
  ignition
- |
  ignobility
- |
  ignoble
- |
  ignobleness
- |
  ignobly
- |
  ignominious
- |
  ignominy
- |
  ignorable
- |
  ignoramus
- |
  ignorance
- |
  ignorant
- |
  ignorantly
- |
  ignore
- |
  ignorer
- |
  Iguacu
- |
  iguana
- |
  Iguazu
- |
  IJssel
- |
  Ijssel
- |
  IJsselmeer
- |
  Ijsselmeer
- |
  Ikhnaton
- |
  ileac
- |
  ileal
- |
  ileitis
- |
  Ilene
- |
  ileum
- |
  iliac
- |
  Iliad
- |
  Ilion
- |
  Ilium
- |
  ilium
- |
  Illampu
- |
  illegal
- |
  illegality
- |
  illegally
- |
  illegibility
- |
  illegible
- |
  illegibly
- |
  illegitimacy
- |
  illegitimate
- |
  illiberal
- |
  illiberality
- |
  illiberally
- |
  illicit
- |
  illicitly
- |
  illicitness
- |
  illimitable
- |
  illimitably
- |
  Illinoian
- |
  Illinois
- |
  Illinoisan
- |
  illiquid
- |
  illiteracy
- |
  illiterate
- |
  illiterately
- |
  illness
- |
  illocution
- |
  illogical
- |
  illogicality
- |
  illogically
- |
  illuminable
- |
  illuminate
- |
  illuminated
- |
  Illuminati
- |
  illuminati
- |
  illuminating
- |
  illumination
- |
  illuminator
- |
  illumine
- |
  illuminism
- |
  illuminist
- |
  illusion
- |
  illusional
- |
  illusionary
- |
  illusionism
- |
  illusionist
- |
  illusive
- |
  illusively
- |
  illusiveness
- |
  illusorily
- |
  illusoriness
- |
  illusory
- |
  illustrate
- |
  illustrated
- |
  illustration
- |
  illustrative
- |
  illustrator
- |
  illustrious
- |
  Illyria
- |
  Illyrian
- |
  image
- |
  imagery
- |
  imaginable
- |
  imaginably
- |
  imaginal
- |
  imaginary
- |
  imagination
- |
  imaginative
- |
  imagine
- |
  imagines
- |
  imaging
- |
  imagism
- |
  imagist
- |
  imagistic
- |
  imago
- |
  imamate
- |
  imbalance
- |
  imbalanced
- |
  imbecile
- |
  imbecilic
- |
  imbecility
- |
  imbed
- |
  imbibe
- |
  imbiber
- |
  imbibition
- |
  imbricate
- |
  imbricated
- |
  imbricating
- |
  imbrication
- |
  imbroglio
- |
  imbrue
- |
  imbue
- |
  imbued
- |
  imitable
- |
  imitate
- |
  imitation
- |
  imitative
- |
  imitatively
- |
  imitator
- |
  immaculacy
- |
  immaculate
- |
  immaculately
- |
  immanence
- |
  immanency
- |
  immanent
- |
  immanentism
- |
  immanentist
- |
  immanently
- |
  Immanuel
- |
  immaterial
- |
  immaterially
- |
  immature
- |
  immaturely
- |
  immaturity
- |
  immeasurable
- |
  immeasurably
- |
  immediacies
- |
  immediacy
- |
  immediate
- |
  immediately
- |
  immemorial
- |
  immemorially
- |
  immense
- |
  immensely
- |
  immenseness
- |
  immensity
- |
  immerse
- |
  immersed
- |
  immersible
- |
  immersion
- |
  immesh
- |
  immigrant
- |
  immigrate
- |
  immigration
- |
  imminence
- |
  imminent
- |
  imminently
- |
  immiscible
- |
  immobile
- |
  immobility
- |
  immobilize
- |
  immoderacy
- |
  immoderate
- |
  immoderately
- |
  immoderation
- |
  immodest
- |
  immodestly
- |
  immodesty
- |
  immolate
- |
  immolation
- |
  immolator
- |
  immoral
- |
  immorality
- |
  immorally
- |
  immortal
- |
  immortality
- |
  immortalize
- |
  immortally
- |
  immovability
- |
  immovable
- |
  immovably
- |
  immune
- |
  immunise
- |
  immunity
- |
  immunization
- |
  immunize
- |
  immunologic
- |
  immunologist
- |
  immunology
- |
  immuration
- |
  immure
- |
  immurement
- |
  immutability
- |
  immutable
- |
  immutably
- |
  Imogen
- |
  impact
- |
  impacted
- |
  impaction
- |
  impair
- |
  impaired
- |
  impairment
- |
  impala
- |
  impale
- |
  impaled
- |
  impalement
- |
  impaler
- |
  impalpable
- |
  impalpably
- |
  impanel
- |
  impanelment
- |
  impart
- |
  impartial
- |
  impartiality
- |
  impartially
- |
  impassable
- |
  impassably
- |
  impasse
- |
  impassible
- |
  impassibly
- |
  impassioned
- |
  impassive
- |
  impassively
- |
  impassivity
- |
  impasto
- |
  impatience
- |
  impatiens
- |
  impatient
- |
  impatiently
- |
  impeach
- |
  impeachable
- |
  impeacher
- |
  impeachment
- |
  impeccable
- |
  impeccably
- |
  impecunious
- |
  impedance
- |
  impede
- |
  impeder
- |
  impediment
- |
  impedimenta
- |
  impedimental
- |
  impel
- |
  impeller
- |
  impellor
- |
  impend
- |
  impending
- |
  impenetrable
- |
  impenetrably
- |
  impenitence
- |
  impenitent
- |
  impenitently
- |
  imperatival
- |
  imperative
- |
  imperatively
- |
  imperceptive
- |
  imperfect
- |
  imperfection
- |
  imperfectly
- |
  imperial
- |
  imperialism
- |
  imperialist
- |
  imperially
- |
  imperialness
- |
  imperil
- |
  imperilment
- |
  imperious
- |
  imperiously
- |
  imperishable
- |
  imperishably
- |
  impermanence
- |
  impermanency
- |
  impermanent
- |
  impermeable
- |
  impermeably
- |
  impersonal
- |
  impersonally
- |
  impersonate
- |
  impersonator
- |
  impertinence
- |
  impertinent
- |
  impervious
- |
  imperviously
- |
  impetigo
- |
  impetuosity
- |
  impetuous
- |
  impetuously
- |
  impetus
- |
  impiety
- |
  impinge
- |
  impingement
- |
  impinger
- |
  impious
- |
  impiously
- |
  impiousness
- |
  impish
- |
  impishly
- |
  impishness
- |
  implacable
- |
  implacably
- |
  implant
- |
  implantable
- |
  implantation
- |
  implausible
- |
  implausibly
- |
  implement
- |
  implicate
- |
  implicated
- |
  implication
- |
  implicative
- |
  implicit
- |
  implicitly
- |
  implicitness
- |
  implode
- |
  implore
- |
  imploringly
- |
  implosion
- |
  implosive
- |
  imply
- |
  impolite
- |
  impolitely
- |
  impoliteness
- |
  impolitic
- |
  impoliticly
- |
  imponderable
- |
  imponderably
- |
  import
- |
  importable
- |
  importance
- |
  important
- |
  importantly
- |
  importation
- |
  importer
- |
  importunate
- |
  importune
- |
  importunely
- |
  importuner
- |
  importunity
- |
  impose
- |
  imposer
- |
  imposing
- |
  imposingly
- |
  imposition
- |
  impossible
- |
  impossibly
- |
  impost
- |
  imposter
- |
  impostor
- |
  imposture
- |
  impotence
- |
  impotency
- |
  impotent
- |
  impotently
- |
  impound
- |
  impoundable
- |
  impoundage
- |
  impounder
- |
  impoundment
- |
  impoverish
- |
  impoverished
- |
  impractical
- |
  imprecate
- |
  imprecation
- |
  imprecator
- |
  imprecatory
- |
  imprecise
- |
  imprecisely
- |
  imprecision
- |
  impregnable
- |
  impregnably
- |
  impregnate
- |
  impregnation
- |
  impregnator
- |
  impresario
- |
  impress
- |
  impressed
- |
  impresser
- |
  impressible
- |
  impression
- |
  impressive
- |
  impressively
- |
  impressment
- |
  imprimatur
- |
  imprint
- |
  imprinter
- |
  imprison
- |
  imprisonable
- |
  imprisonment
- |
  improbable
- |
  improbably
- |
  impromptu
- |
  improper
- |
  improperly
- |
  improperness
- |
  impropriety
- |
  improvable
- |
  improve
- |
  improved
- |
  improvement
- |
  improvidence
- |
  improvident
- |
  improvise
- |
  improviser
- |
  improvisor
- |
  imprudence
- |
  imprudent
- |
  imprudently
- |
  impudence
- |
  impudent
- |
  impudently
- |
  impugn
- |
  impugnable
- |
  impugner
- |
  impugnment
- |
  impuissance
- |
  impulse
- |
  impulsion
- |
  impulsive
- |
  impulsively
- |
  impulsivity
- |
  impunity
- |
  impure
- |
  impurely
- |
  impureness
- |
  impurity
- |
  imputable
- |
  imputation
- |
  impute
- |
  inability
- |
  inaccessible
- |
  inaccessibly
- |
  inaccuracy
- |
  inaccurate
- |
  inaccurately
- |
  inaction
- |
  inactivate
- |
  inactivation
- |
  inactive
- |
  inactively
- |
  inactiveness
- |
  inactivity
- |
  inadequacy
- |
  inadequate
- |
  inadequately
- |
  inadmissible
- |
  inadmissibly
- |
  inadvertence
- |
  inadvertency
- |
  inadvertent
- |
  inadvisable
- |
  inalienable
- |
  inalienably
- |
  inamorata
- |
  inamorato
- |
  inane
- |
  inanely
- |
  inaneness
- |
  inanimate
- |
  inanimately
- |
  inanition
- |
  inanity
- |
  inapparent
- |
  inapplicable
- |
  inapposite
- |
  inapt
- |
  inaptitude
- |
  inaptly
- |
  inaptness
- |
  inarguable
- |
  inarticulacy
- |
  inarticulate
- |
  inartistic
- |
  inattention
- |
  inattentive
- |
  inaudibility
- |
  inaudible
- |
  inaudibly
- |
  inaugural
- |
  inaugurate
- |
  inauguration
- |
  inaugurator
- |
  inauspicious
- |
  inauthentic
- |
  inboard
- |
  inborn
- |
  inbound
- |
  inbred
- |
  inbreed
- |
  inbreeder
- |
  inbreeding
- |
  incalculable
- |
  incalculably
- |
  Incan
- |
  incandescent
- |
  incantation
- |
  incantatory
- |
  incapability
- |
  incapable
- |
  incapably
- |
  incapacitant
- |
  incapacitate
- |
  incapacity
- |
  incarcerate
- |
  incarcerator
- |
  incarnadine
- |
  incarnate
- |
  Incarnation
- |
  incarnation
- |
  incase
- |
  incautious
- |
  incautiously
- |
  incendiarism
- |
  incendiary
- |
  incense
- |
  incensed
- |
  incentive
- |
  incentivize
- |
  inception
- |
  inceptive
- |
  incertitude
- |
  incessance
- |
  incessancy
- |
  incessant
- |
  incessantly
- |
  incest
- |
  incestuous
- |
  incestuously
- |
  inchoate
- |
  inchoately
- |
  inchoateness
- |
  Inchon
- |
  inchworm
- |
  incidence
- |
  incident
- |
  incidental
- |
  incidentally
- |
  incidentals
- |
  incinerate
- |
  incineration
- |
  incinerator
- |
  incipience
- |
  incipiency
- |
  incipient
- |
  incipiently
- |
  incise
- |
  incision
- |
  incisive
- |
  incisively
- |
  incisiveness
- |
  incisor
- |
  incitation
- |
  incite
- |
  incitement
- |
  inciter
- |
  incivilities
- |
  incivility
- |
  inclemency
- |
  inclement
- |
  inclemently
- |
  inclination
- |
  incline
- |
  inclined
- |
  incliner
- |
  inclose
- |
  inclosure
- |
  include
- |
  included
- |
  including
- |
  inclusion
- |
  inclusive
- |
  inclusively
- |
  incognito
- |
  incoherence
- |
  incoherency
- |
  incoherent
- |
  incoherently
- |
  income
- |
  incoming
- |
  incommode
- |
  incommodious
- |
  incomparable
- |
  incomparably
- |
  incompatible
- |
  incompatibly
- |
  incompetence
- |
  incompetency
- |
  incompetent
- |
  incomplete
- |
  incompletely
- |
  incompletion
- |
  inconclusive
- |
  incongruence
- |
  incongruent
- |
  incongruity
- |
  incongruous
- |
  inconsistent
- |
  inconsolable
- |
  inconsolably
- |
  inconstancy
- |
  inconstant
- |
  inconstantly
- |
  incontinence
- |
  incontinent
- |
  inconvenient
- |
  incorporate
- |
  Incorporated
- |
  incorporated
- |
  incorporator
- |
  incorporeal
- |
  incorporeity
- |
  incorrect
- |
  incorrectly
- |
  incorrigible
- |
  incorrigibly
- |
  increase
- |
  increased
- |
  increasing
- |
  increasingly
- |
  incredible
- |
  incredibly
- |
  incredulity
- |
  incredulous
- |
  increment
- |
  incremental
- |
  incriminate
- |
  incrust
- |
  incrustation
- |
  incubate
- |
  incubation
- |
  incubative
- |
  incubator
- |
  incubi
- |
  incubus
- |
  incudes
- |
  inculcate
- |
  inculcation
- |
  inculcative
- |
  inculcator
- |
  inculpable
- |
  inculpate
- |
  inculpation
- |
  inculpatory
- |
  incumbency
- |
  incumbent
- |
  incumber
- |
  incumbrance
- |
  incunabula
- |
  incunabulum
- |
  incur
- |
  incurability
- |
  incurable
- |
  incurably
- |
  incurious
- |
  incuriously
- |
  incursion
- |
  incus
- |
  indebted
- |
  indebtedness
- |
  indecency
- |
  indecent
- |
  indecently
- |
  indecision
- |
  indecisive
- |
  indecisively
- |
  indecorous
- |
  indecorously
- |
  indeed
- |
  indefeasible
- |
  indefeasibly
- |
  indefensible
- |
  indefensibly
- |
  indefinable
- |
  indefinably
- |
  indefinite
- |
  indefinitely
- |
  indelibility
- |
  indelible
- |
  indelibly
- |
  indelicacy
- |
  indelicate
- |
  indelicately
- |
  indemnifier
- |
  indemnify
- |
  indemnity
- |
  indent
- |
  indentation
- |
  indention
- |
  indenture
- |
  Independence
- |
  independence
- |
  independent
- |
  index
- |
  indexation
- |
  indexer
- |
  indexing
- |
  India
- |
  Indian
- |
  Indiana
- |
  Indianan
- |
  Indianapolis
- |
  Indianian
- |
  Indianize
- |
  Indianness
- |
  Indic
- |
  indicate
- |
  indication
- |
  indicative
- |
  indicatively
- |
  indicator
- |
  indices
- |
  indicia
- |
  indict
- |
  indictable
- |
  indictee
- |
  indicter
- |
  indictment
- |
  indictor
- |
  indie
- |
  Indies
- |
  indifference
- |
  indifferent
- |
  indigence
- |
  indigenous
- |
  indigenously
- |
  indigent
- |
  indigently
- |
  indigestible
- |
  indigestibly
- |
  indigestion
- |
  indignant
- |
  indignantly
- |
  indignation
- |
  indignity
- |
  indigo
- |
  indirect
- |
  indirection
- |
  indirectly
- |
  indirectness
- |
  indiscreet
- |
  indiscreetly
- |
  indiscretion
- |
  indisposed
- |
  indisputable
- |
  indisputably
- |
  indissoluble
- |
  indissolubly
- |
  indistinct
- |
  indistinctly
- |
  indite
- |
  indium
- |
  individual
- |
  individually
- |
  individuate
- |
  indivisible
- |
  indivisibly
- |
  Indochina
- |
  Indochinese
- |
  indoctrinate
- |
  indolence
- |
  indolent
- |
  indolently
- |
  indomitable
- |
  indomitably
- |
  Indonesia
- |
  Indonesian
- |
  indoor
- |
  indoors
- |
  Indore
- |
  indorse
- |
  indubitable
- |
  indubitably
- |
  induce
- |
  induced
- |
  inducement
- |
  inducer
- |
  inducible
- |
  induct
- |
  inductance
- |
  inductee
- |
  induction
- |
  inductive
- |
  inductively
- |
  inductor
- |
  indue
- |
  indulge
- |
  indulgence
- |
  indulgent
- |
  indulgently
- |
  indulger
- |
  indurate
- |
  indurated
- |
  induration
- |
  indurative
- |
  Indus
- |
  industrial
- |
  industrially
- |
  industrious
- |
  industry
- |
  indwell
- |
  inebriate
- |
  inebriated
- |
  inebriation
- |
  inebriety
- |
  inedibility
- |
  inedible
- |
  inedibly
- |
  ineducable
- |
  ineffability
- |
  ineffable
- |
  ineffably
- |
  ineffaceable
- |
  ineffective
- |
  ineffectual
- |
  inefficacy
- |
  inefficiency
- |
  inefficient
- |
  inelastic
- |
  inelasticity
- |
  inelegance
- |
  inelegant
- |
  inelegantly
- |
  ineligible
- |
  ineligibly
- |
  ineluctable
- |
  ineluctably
- |
  inept
- |
  ineptitude
- |
  ineptly
- |
  ineptness
- |
  inequality
- |
  inequitable
- |
  inequitably
- |
  inequity
- |
  ineradicable
- |
  inerrancy
- |
  inerrant
- |
  inert
- |
  inertia
- |
  inertial
- |
  inertialess
- |
  inertly
- |
  inertness
- |
  inescapable
- |
  inescapably
- |
  inessential
- |
  inestimable
- |
  inestimably
- |
  inevitable
- |
  inevitably
- |
  inexact
- |
  inexactly
- |
  inexactness
- |
  inexcusable
- |
  inexcusably
- |
  inexorable
- |
  inexorably
- |
  inexpedience
- |
  inexpediency
- |
  inexpedient
- |
  inexpensive
- |
  inexperience
- |
  inexpert
- |
  inexpertly
- |
  inexpiable
- |
  inexplicable
- |
  inexplicably
- |
  inexpressive
- |
  inextricable
- |
  inextricably
- |
  infallible
- |
  infallibly
- |
  infamous
- |
  infamously
- |
  infamousness
- |
  infamy
- |
  infancy
- |
  infant
- |
  infanticide
- |
  infantile
- |
  infantilism
- |
  infantry
- |
  infantryman
- |
  infarct
- |
  infarcted
- |
  infarction
- |
  infatuate
- |
  infatuated
- |
  infatuation
- |
  infeasible
- |
  infect
- |
  infected
- |
  infection
- |
  infectious
- |
  infectiously
- |
  infective
- |
  infelicitous
- |
  infelicity
- |
  infer
- |
  inferable
- |
  inference
- |
  inferential
- |
  inferior
- |
  inferiority
- |
  infernal
- |
  infernally
- |
  inferno
- |
  inferrable
- |
  infertile
- |
  infertility
- |
  infest
- |
  infestation
- |
  infested
- |
  infester
- |
  infidel
- |
  infidelity
- |
  infield
- |
  infielder
- |
  infighter
- |
  infighting
- |
  infiltrate
- |
  infiltration
- |
  infiltrator
- |
  infinite
- |
  infinitely
- |
  infiniteness
- |
  infinitival
- |
  infinitive
- |
  infinitude
- |
  infinity
- |
  infirm
- |
  infirmary
- |
  infirmity
- |
  infirmly
- |
  infirmness
- |
  inflame
- |
  inflamed
- |
  inflammable
- |
  inflammably
- |
  inflammation
- |
  inflammatory
- |
  inflatable
- |
  inflate
- |
  inflated
- |
  inflater
- |
  inflation
- |
  inflationary
- |
  inflationism
- |
  inflationist
- |
  inflator
- |
  inflect
- |
  inflection
- |
  inflectional
- |
  inflective
- |
  inflexible
- |
  inflexibly
- |
  inflexion
- |
  inflict
- |
  inflicter
- |
  infliction
- |
  inflictive
- |
  inflictor
- |
  inflight
- |
  inflorescent
- |
  inflow
- |
  influence
- |
  influential
- |
  influenza
- |
  influx
- |
  infold
- |
  infomercial
- |
  inform
- |
  informal
- |
  informality
- |
  informally
- |
  informant
- |
  information
- |
  informative
- |
  informed
- |
  informer
- |
  infotainment
- |
  infra
- |
  infraction
- |
  infractor
- |
  infrangible
- |
  infrangibly
- |
  infrared
- |
  infrasonic
- |
  infrequence
- |
  infrequency
- |
  infrequent
- |
  infrequently
- |
  infringe
- |
  infringement
- |
  infringer
- |
  infuriate
- |
  infuriated
- |
  infuriating
- |
  infuse
- |
  infuser
- |
  infusible
- |
  infusion
- |
  ingather
- |
  ingenious
- |
  ingeniously
- |
  ingenue
- |
  ingenuity
- |
  ingenuous
- |
  ingenuously
- |
  ingest
- |
  ingestion
- |
  inglenook
- |
  Inglewood
- |
  inglorious
- |
  ingloriously
- |
  ingot
- |
  ingrain
- |
  ingrained
- |
  ingrate
- |
  ingratiate
- |
  ingratiating
- |
  ingratiation
- |
  ingratiatory
- |
  ingratitude
- |
  ingredient
- |
  Ingres
- |
  ingress
- |
  ingression
- |
  Ingrid
- |
  ingrowing
- |
  ingrown
- |
  inguinal
- |
  inhabit
- |
  inhabitable
- |
  inhabitant
- |
  inhalant
- |
  inhalation
- |
  inhalator
- |
  inhale
- |
  inhaler
- |
  inharmonious
- |
  inhere
- |
  inherence
- |
  inherency
- |
  inherent
- |
  inherently
- |
  inherit
- |
  inheritable
- |
  inheritance
- |
  inheritor
- |
  inhibit
- |
  inhibited
- |
  inhibiter
- |
  inhibition
- |
  inhibitive
- |
  inhibitor
- |
  inhibitory
- |
  inhospitable
- |
  inhospitably
- |
  inhuman
- |
  inhumane
- |
  inhumanely
- |
  inhumanity
- |
  inhumanly
- |
  inhumanness
- |
  inimical
- |
  inimically
- |
  inimitable
- |
  inimitably
- |
  iniquitous
- |
  iniquitously
- |
  iniquity
- |
  initial
- |
  initialize
- |
  initially
- |
  initiate
- |
  initiation
- |
  initiative
- |
  initiator
- |
  initiatory
- |
  inject
- |
  injection
- |
  injector
- |
  injudicious
- |
  injunction
- |
  injunctive
- |
  injure
- |
  injured
- |
  injurer
- |
  injurious
- |
  injuriously
- |
  injury
- |
  injustice
- |
  inkblot
- |
  inkhorn
- |
  inkiness
- |
  inkling
- |
  inkstand
- |
  inkwell
- |
  inlaid
- |
  Inland
- |
  inland
- |
  inlay
- |
  inlet
- |
  inmate
- |
  inmost
- |
  innards
- |
  innate
- |
  innately
- |
  innateness
- |
  inner
- |
  innermost
- |
  innerness
- |
  innersole
- |
  innerspring
- |
  innervate
- |
  innervation
- |
  inning
- |
  innings
- |
  innkeeper
- |
  innocence
- |
  Innocent
- |
  innocent
- |
  innocently
- |
  innocuous
- |
  innocuously
- |
  innominate
- |
  innovate
- |
  innovation
- |
  innovational
- |
  innovative
- |
  innovator
- |
  Innsbruck
- |
  innuendo
- |
  innumerable
- |
  innumerably
- |
  innumeracy
- |
  innumerate
- |
  inocula
- |
  inoculable
- |
  inoculant
- |
  inoculate
- |
  inoculation
- |
  inoculator
- |
  inoculum
- |
  inoffensive
- |
  inoperable
- |
  inoperative
- |
  inopportune
- |
  inordinate
- |
  inordinately
- |
  inorganic
- |
  inpatient
- |
  input
- |
  inquest
- |
  inquietude
- |
  inquire
- |
  inquirer
- |
  inquiring
- |
  inquiringly
- |
  inquiry
- |
  Inquisition
- |
  inquisition
- |
  inquisitive
- |
  inquisitor
- |
  inroad
- |
  inroads
- |
  inrush
- |
  insalubrious
- |
  insane
- |
  insanely
- |
  insanitary
- |
  insanity
- |
  insatiable
- |
  insatiably
- |
  insatiate
- |
  insatiately
- |
  insatiety
- |
  inscribe
- |
  inscriber
- |
  inscription
- |
  inscrutable
- |
  inscrutably
- |
  inseam
- |
  insect
- |
  insecticidal
- |
  insecticide
- |
  insectivore
- |
  insecure
- |
  insecurely
- |
  insecurity
- |
  inseminate
- |
  insemination
- |
  inseminator
- |
  insensate
- |
  insensately
- |
  insensible
- |
  insensibly
- |
  insensitive
- |
  insentience
- |
  insentient
- |
  inseparable
- |
  inseparably
- |
  insert
- |
  insertion
- |
  inset
- |
  inshore
- |
  inside
- |
  insider
- |
  insides
- |
  insidious
- |
  insidiously
- |
  insight
- |
  insightful
- |
  insigne
- |
  insignia
- |
  insincere
- |
  insincerely
- |
  insincerity
- |
  insinuate
- |
  insinuating
- |
  insinuation
- |
  insinuative
- |
  insinuator
- |
  insipid
- |
  insipidity
- |
  insipidly
- |
  insipidness
- |
  insist
- |
  insistence
- |
  insistency
- |
  insistent
- |
  insistently
- |
  insistingly
- |
  insobriety
- |
  insofar
- |
  insolation
- |
  insole
- |
  insolence
- |
  insolent
- |
  insolently
- |
  insolubility
- |
  insolubilize
- |
  insoluble
- |
  insolubly
- |
  insolvable
- |
  insolvency
- |
  insolvent
- |
  insomnia
- |
  insomniac
- |
  insomuch
- |
  insouciance
- |
  insouciant
- |
  insouciantly
- |
  inspect
- |
  inspection
- |
  inspector
- |
  inspectorate
- |
  inspiration
- |
  inspire
- |
  inspired
- |
  inspirer
- |
  inspiring
- |
  inspirit
- |
  instability
- |
  instal
- |
  install
- |
  installation
- |
  installer
- |
  installment
- |
  instalment
- |
  instance
- |
  instant
- |
  instanter
- |
  instantiate
- |
  instantly
- |
  instate
- |
  instatement
- |
  instead
- |
  instep
- |
  instigate
- |
  instigation
- |
  instigator
- |
  instil
- |
  instill
- |
  instillation
- |
  instiller
- |
  instillment
- |
  instinct
- |
  instinctive
- |
  instinctual
- |
  institute
- |
  instituter
- |
  institutes
- |
  institution
- |
  institutor
- |
  instruct
- |
  instruction
- |
  instructions
- |
  instructive
- |
  instructor
- |
  instrument
- |
  instrumental
- |
  insufferable
- |
  insufferably
- |
  insufficient
- |
  insufflate
- |
  insufflation
- |
  insular
- |
  insularity
- |
  insularly
- |
  insulate
- |
  insulation
- |
  insulator
- |
  insulin
- |
  insult
- |
  insulted
- |
  insulting
- |
  insultingly
- |
  insuperable
- |
  insuperably
- |
  insurability
- |
  insurable
- |
  insurance
- |
  insure
- |
  insured
- |
  insurer
- |
  insurgence
- |
  insurgency
- |
  insurgent
- |
  insurgents
- |
  insurrection
- |
  intact
- |
  intactness
- |
  intaglio
- |
  intaglioed
- |
  intake
- |
  intangible
- |
  intangibly
- |
  intarsia
- |
  integer
- |
  integrable
- |
  integral
- |
  integrality
- |
  integrally
- |
  integrate
- |
  integrated
- |
  integration
- |
  integrative
- |
  integrity
- |
  integument
- |
  integumental
- |
  intellect
- |
  intellection
- |
  intellective
- |
  intellectual
- |
  intelligence
- |
  intelligent
- |
  intelligible
- |
  intelligibly
- |
  intemperance
- |
  intemperate
- |
  intend
- |
  intendant
- |
  intended
- |
  intense
- |
  intensely
- |
  intenseness
- |
  intensifier
- |
  intensify
- |
  intension
- |
  intensional
- |
  intensity
- |
  intensive
- |
  intensively
- |
  intent
- |
  intention
- |
  intentional
- |
  intentions
- |
  intently
- |
  intentness
- |
  inter
- |
  interact
- |
  interaction
- |
  interactive
- |
  interatomic
- |
  interbred
- |
  interbreed
- |
  intercalary
- |
  intercalate
- |
  intercede
- |
  interceder
- |
  intercept
- |
  interception
- |
  interceptive
- |
  interceptor
- |
  intercession
- |
  intercessor
- |
  intercessory
- |
  interchange
- |
  intercom
- |
  interconnect
- |
  intercostal
- |
  intercourse
- |
  interdict
- |
  interdiction
- |
  interdictory
- |
  interest
- |
  interested
- |
  interesting
- |
  interests
- |
  interface
- |
  interfacial
- |
  interfaith
- |
  interfere
- |
  interference
- |
  interferer
- |
  interferon
- |
  interfile
- |
  interfuse
- |
  interfusion
- |
  interglacial
- |
  interim
- |
  interior
- |
  interiorize
- |
  interject
- |
  interjection
- |
  interjectory
- |
  interlace
- |
  interlaced
- |
  interlard
- |
  interleave
- |
  interleaving
- |
  interleukin
- |
  interline
- |
  interlinear
- |
  interlining
- |
  interlink
- |
  interlock
- |
  interlocking
- |
  interlocutor
- |
  interlope
- |
  interloper
- |
  interlude
- |
  intermarry
- |
  intermediary
- |
  intermediate
- |
  interment
- |
  intermezzi
- |
  intermezzo
- |
  interminable
- |
  interminably
- |
  intermingle
- |
  intermission
- |
  intermit
- |
  intermittent
- |
  intermix
- |
  intermixture
- |
  intermontane
- |
  intern
- |
  internal
- |
  internalize
- |
  internally
- |
  interne
- |
  internecine
- |
  internee
- |
  Internet
- |
  internist
- |
  internment
- |
  internship
- |
  internuncio
- |
  interoffice
- |
  interplay
- |
  Interpol
- |
  interpolate
- |
  interpolator
- |
  interposable
- |
  interpose
- |
  interposer
- |
  interpret
- |
  interpreter
- |
  interpretive
- |
  interrace
- |
  interracial
- |
  interregna
- |
  interregnal
- |
  interregnum
- |
  interrelate
- |
  interrelated
- |
  interrogate
- |
  interrogator
- |
  interrupt
- |
  interrupter
- |
  interruption
- |
  interruptive
- |
  intersect
- |
  intersection
- |
  interservice
- |
  intersession
- |
  intersperse
- |
  interspersed
- |
  interstate
- |
  interstellar
- |
  interstice
- |
  interstices
- |
  interstitial
- |
  intertidal
- |
  intertwine
- |
  intertwined
- |
  intertwist
- |
  interurban
- |
  interval
- |
  intervallic
- |
  intervene
- |
  intervener
- |
  intervenient
- |
  intervening
- |
  intervenor
- |
  intervention
- |
  interview
- |
  interviewee
- |
  interviewer
- |
  intervocalic
- |
  interweave
- |
  interwove
- |
  interwoven
- |
  intestacy
- |
  intestate
- |
  intestinal
- |
  intestinally
- |
  intestine
- |
  intestines
- |
  intifada
- |
  intimacy
- |
  intimate
- |
  intimately
- |
  intimation
- |
  intimidate
- |
  intimidated
- |
  intimidating
- |
  intimidation
- |
  intimidator
- |
  intimidatory
- |
  intolerable
- |
  intolerably
- |
  intolerance
- |
  intolerant
- |
  intolerantly
- |
  intonation
- |
  intonational
- |
  intone
- |
  intoner
- |
  intoxicant
- |
  intoxicate
- |
  intoxicated
- |
  intoxicating
- |
  intoxication
- |
  intracity
- |
  intractable
- |
  intractably
- |
  intradermal
- |
  intramural
- |
  intranet
- |
  intransigent
- |
  intransitive
- |
  intraocular
- |
  intrapreneur
- |
  intrastate
- |
  intrauterine
- |
  intravenous
- |
  intrench
- |
  intrepid
- |
  intrepidity
- |
  intrepidly
- |
  intrepidness
- |
  intricacy
- |
  intricate
- |
  intricately
- |
  intrigue
- |
  intrigued
- |
  intriguer
- |
  intriguing
- |
  intriguingly
- |
  intrinsic
- |
  intro
- |
  introduce
- |
  introducible
- |
  introduction
- |
  introductory
- |
  introit
- |
  introject
- |
  introjection
- |
  intromission
- |
  introspect
- |
  introversion
- |
  introversive
- |
  introvert
- |
  introverted
- |
  intrude
- |
  intruder
- |
  intrusion
- |
  intrusive
- |
  intrusively
- |
  intrust
- |
  intubate
- |
  intuit
- |
  intuitable
- |
  intuition
- |
  intuitional
- |
  intuitive
- |
  intuitively
- |
  intumesce
- |
  intumescence
- |
  intumescent
- |
  Inuit
- |
  Inuktitut
- |
  inundate
- |
  inundation
- |
  Inupiaq
- |
  inure
- |
  inurement
- |
  invade
- |
  invader
- |
  invalid
- |
  invalidate
- |
  invalidation
- |
  invalidator
- |
  invalidism
- |
  invalidity
- |
  invalidly
- |
  invaluable
- |
  invaluably
- |
  invariable
- |
  invariably
- |
  invasion
- |
  invasive
- |
  invective
- |
  inveigh
- |
  inveigle
- |
  inveiglement
- |
  inveigler
- |
  invent
- |
  invention
- |
  inventive
- |
  inventively
- |
  inventor
- |
  inventory
- |
  Inverness
- |
  inverse
- |
  inversely
- |
  inversion
- |
  invert
- |
  invertebrate
- |
  inverter
- |
  invertible
- |
  invest
- |
  investigate
- |
  investigator
- |
  investiture
- |
  investment
- |
  investor
- |
  inveteracy
- |
  inveterate
- |
  inveterately
- |
  invidious
- |
  invidiously
- |
  invigorate
- |
  invigorated
- |
  invigorating
- |
  invigoration
- |
  invigorative
- |
  invincible
- |
  invincibly
- |
  inviolable
- |
  inviolably
- |
  inviolacy
- |
  inviolate
- |
  inviolately
- |
  invisibility
- |
  invisible
- |
  invisibly
- |
  invitation
- |
  invitational
- |
  invite
- |
  invitee
- |
  inviting
- |
  invitingly
- |
  invocation
- |
  invocative
- |
  invocatory
- |
  invoice
- |
  invoke
- |
  invoker
- |
  involuntary
- |
  involute
- |
  involution
- |
  involutional
- |
  involve
- |
  involved
- |
  involvement
- |
  invulnerable
- |
  invulnerably
- |
  inward
- |
  inwardly
- |
  inwards
- |
  iodide
- |
  iodine
- |
  iodize
- |
  Ionesco
- |
  Ionia
- |
  Ionian
- |
  Ionic
- |
  ionic
- |
  ionizable
- |
  ionization
- |
  ionize
- |
  ionizer
- |
  ionosphere
- |
  ionospheric
- |
  Iowan
- |
  ipecac
- |
  Iphigenia
- |
  Ipswich
- |
  Iqaluit
- |
  Iquitos
- |
  Iraklion
- |
  Irani
- |
  Iranian
- |
  Iraqi
- |
  irascibility
- |
  irascible
- |
  irascibly
- |
  irate
- |
  irately
- |
  irateness
- |
  Irbid
- |
  Irbil
- |
  ireful
- |
  irefully
- |
  Ireland
- |
  Irene
- |
  irenic
- |
  irenical
- |
  irenically
- |
  irenicism
- |
  irenics
- |
  irides
- |
  iridescence
- |
  iridescent
- |
  iridescently
- |
  iridium
- |
  Irish
- |
  Irishman
- |
  Irishwoman
- |
  irksome
- |
  irksomely
- |
  irksomeness
- |
  Irkutsk
- |
  ironclad
- |
  ironer
- |
  ironic
- |
  ironical
- |
  ironically
- |
  ironicalness
- |
  ironing
- |
  ironist
- |
  irons
- |
  ironstone
- |
  ironware
- |
  ironweed
- |
  ironwood
- |
  ironwork
- |
  ironworker
- |
  ironworks
- |
  irony
- |
  Iroquoian
- |
  Iroquois
- |
  irradiate
- |
  irradiation
- |
  irradiative
- |
  irradiator
- |
  irrational
- |
  irrationally
- |
  Irrawaddy
- |
  irredeemable
- |
  irredeemably
- |
  irredentism
- |
  irredentist
- |
  irreducible
- |
  irreducibly
- |
  irrefragable
- |
  irrefragably
- |
  irrefutable
- |
  irrefutably
- |
  irregardless
- |
  irregular
- |
  irregularity
- |
  irregularly
- |
  irregulars
- |
  irrelevance
- |
  irrelevancy
- |
  irrelevant
- |
  irrelevantly
- |
  irreligion
- |
  irreligious
- |
  irremediable
- |
  irremediably
- |
  irremovable
- |
  irreparable
- |
  irreparably
- |
  irresistible
- |
  irresistibly
- |
  irresolute
- |
  irresolutely
- |
  irresolution
- |
  irrespective
- |
  irreverence
- |
  irreverent
- |
  irreverently
- |
  irreversible
- |
  irreversibly
- |
  irrevocable
- |
  irrevocably
- |
  irrigable
- |
  irrigate
- |
  irrigation
- |
  irrigational
- |
  irrigator
- |
  irritability
- |
  irritable
- |
  irritably
- |
  irritant
- |
  irritate
- |
  irritated
- |
  irritating
- |
  irritatingly
- |
  irritation
- |
  irritative
- |
  irritator
- |
  irrupt
- |
  irruption
- |
  irruptive
- |
  Irtish
- |
  Irtysh
- |
  Irvin
- |
  Irvine
- |
  Irving
- |
  Irwin
- |
  Isaac
- |
  Isabel
- |
  Isabella
- |
  Isabelle
- |
  Isador
- |
  Isadora
- |
  Isadore
- |
  Isaiah
- |
  Isaias
- |
  ischemia
- |
  ischemic
- |
  Iseult
- |
  Isfahan
- |
  Isherwood
- |
  Ishmael
- |
  Ishtar
- |
  Isidor
- |
  isinglass
- |
  Islam
- |
  Islamabad
- |
  Islamic
- |
  island
- |
  islander
- |
  islet
- |
  Islington
- |
  isobar
- |
  isobaric
- |
  isobarism
- |
  isogon
- |
  isogonic
- |
  isolate
- |
  isolated
- |
  isolation
- |
  isolationism
- |
  isolationist
- |
  isolator
- |
  isomer
- |
  isomeric
- |
  isomerism
- |
  isometric
- |
  isometrical
- |
  isometrics
- |
  isomorph
- |
  isomorphic
- |
  isomorphism
- |
  isomorphous
- |
  isoprene
- |
  isosceles
- |
  isostasy
- |
  isostatic
- |
  isotherm
- |
  isothermal
- |
  isotope
- |
  isotopic
- |
  isotopically
- |
  isotopy
- |
  isotropic
- |
  isotropism
- |
  isotropy
- |
  Ispahan
- |
  Israel
- |
  Israeli
- |
  Israelite
- |
  issei
- |
  issuance
- |
  issue
- |
  issuer
- |
  Istanbul
- |
  isthmi
- |
  isthmian
- |
  isthmus
- |
  Istria
- |
  Istrian
- |
  Italian
- |
  Italianate
- |
  Italic
- |
  italic
- |
  italicize
- |
  italicized
- |
  italics
- |
  Italy
- |
  itchiness
- |
  itching
- |
  itchy
- |
  itemization
- |
  itemize
- |
  itemized
- |
  itemizer
- |
  iterate
- |
  iteration
- |
  iterative
- |
  iteratively
- |
  Ithaca
- |
  Ithaki
- |
  itineracy
- |
  itinerancy
- |
  itinerant
- |
  itinerantly
- |
  itinerary
- |
  itself
- |
  Ivanovo
- |
  ivied
- |
  Ivorian
- |
  ivories
- |
  ivory
- |
  Ixtapalapa
- |
  Iyyar
- |
  Izhevsk
- |
  Izmir
- |
  Izmit
- |
  Jabalpur
- |
  jabber
- |
  jabberer
- |
  jabberwocky
- |
  jabot
- |
  jacaranda
- |
  jackal
- |
  jackanapes
- |
  jackass
- |
  jackboot
- |
  jackdaw
- |
  jacket
- |
  jacketed
- |
  jackhammer
- |
  Jackie
- |
  jackknife
- |
  jackknives
- |
  jackleg
- |
  jackpot
- |
  jackrabbit
- |
  jacks
- |
  jackscrew
- |
  Jackson
- |
  Jacksonville
- |
  jackstraw
- |
  Jacky
- |
  Jacob
- |
  Jacobean
- |
  Jacobin
- |
  Jacobinic
- |
  Jacobinical
- |
  Jacobinism
- |
  Jacobite
- |
  Jacobitical
- |
  Jacobitism
- |
  Jacquard
- |
  jacquard
- |
  Jacque
- |
  Jacquelin
- |
  Jacqueline
- |
  Jacquelyn
- |
  Jacques
- |
  Jacuzzi
- |
  jaded
- |
  jadedly
- |
  jadedness
- |
  jadeite
- |
  Jaffa
- |
  jagged
- |
  jaggedly
- |
  jaggedness
- |
  jaggies
- |
  jaguar
- |
  jailbird
- |
  jailbreak
- |
  jailer
- |
  jailor
- |
  Jaipur
- |
  Jakarta
- |
  jalap
- |
  Jalapa
- |
  jalapeno
- |
  Jalisco
- |
  jalopy
- |
  jalousie
- |
  Jamaica
- |
  Jamaican
- |
  jambalaya
- |
  jamboree
- |
  James
- |
  Jamestown
- |
  Jamie
- |
  jammed
- |
  jammer
- |
  jamming
- |
  jampacked
- |
  Jamshedpur
- |
  Janacek
- |
  Janet
- |
  Janette
- |
  jangle
- |
  jangler
- |
  Janice
- |
  Janie
- |
  Janis
- |
  janitor
- |
  janitorial
- |
  January
- |
  Janus
- |
  Japan
- |
  japan
- |
  Japanese
- |
  japanned
- |
  japer
- |
  japery
- |
  jardiniere
- |
  Jared
- |
  jarful
- |
  jargon
- |
  jargonistic
- |
  jargonize
- |
  Jarlsberg
- |
  jarring
- |
  jarringly
- |
  Jarvis
- |
  jasmine
- |
  Jason
- |
  Jasper
- |
  jasper
- |
  jaundice
- |
  jaundiced
- |
  jaunt
- |
  jauntily
- |
  jauntiness
- |
  jaunty
- |
  Javan
- |
  Javanese
- |
  javelin
- |
  jawbone
- |
  jawbreaker
- |
  jawed
- |
  jawless
- |
  jaybird
- |
  Jayne
- |
  jayvee
- |
  jaywalk
- |
  jaywalker
- |
  jaywalking
- |
  jazzed
- |
  jazzily
- |
  jazziness
- |
  jazzy
- |
  jealous
- |
  jealously
- |
  jealousness
- |
  jealousy
- |
  Jeanette
- |
  Jeanie
- |
  Jeanine
- |
  Jeanne
- |
  Jeannette
- |
  Jeannie
- |
  Jeannine
- |
  jeans
- |
  Jedda
- |
  jeerer
- |
  jeering
- |
  jeeringly
- |
  Jeeves
- |
  Jefferson
- |
  Jeffersonian
- |
  Jeffery
- |
  Jeffrey
- |
  Jeffry
- |
  jehad
- |
  Jehosaphat
- |
  Jehovah
- |
  jejuna
- |
  jejunal
- |
  jejune
- |
  jejunely
- |
  jejuneness
- |
  jejunum
- |
  jellabah
- |
  jello
- |
  jelly
- |
  jellybean
- |
  jellyfish
- |
  jellylike
- |
  jellyroll
- |
  Jemima
- |
  jennet
- |
  Jennie
- |
  Jennifer
- |
  Jenny
- |
  jenny
- |
  jeopardise
- |
  jeopardize
- |
  jeopardy
- |
  Jerald
- |
  Jeraldine
- |
  jerboa
- |
  jeremiad
- |
  Jeremiah
- |
  Jeremias
- |
  Jeremy
- |
  Jericho
- |
  Jerilyn
- |
  jerkily
- |
  jerkin
- |
  jerkiness
- |
  jerkwater
- |
  jerky
- |
  jeroboam
- |
  Jerold
- |
  Jerome
- |
  Jerrie
- |
  Jerrold
- |
  Jerry
- |
  jerrybuilt
- |
  Jersey
- |
  jersey
- |
  Jerseyite
- |
  Jerusalem
- |
  Jerusalemite
- |
  Jervis
- |
  Jessamine
- |
  jessamine
- |
  Jesse
- |
  Jessica
- |
  Jessie
- |
  jester
- |
  jestingly
- |
  Jesuit
- |
  Jesus
- |
  jetlag
- |
  jetliner
- |
  jetport
- |
  jetsam
- |
  jettison
- |
  jetty
- |
  Jewel
- |
  jewel
- |
  jeweled
- |
  jeweler
- |
  Jewell
- |
  jeweller
- |
  jewellery
- |
  jewelry
- |
  jewels
- |
  jewelweed
- |
  Jewess
- |
  Jewish
- |
  Jewishness
- |
  Jewry
- |
  Jezebel
- |
  jezebel
- |
  jibber
- |
  jibing
- |
  Jidda
- |
  jiffy
- |
  jigger
- |
  jiggle
- |
  jiggly
- |
  jigsaw
- |
  jihad
- |
  Jilin
- |
  jillion
- |
  Jimmie
- |
  jimmies
- |
  Jimmy
- |
  jimmy
- |
  jimsonweed
- |
  Jinan
- |
  jingle
- |
  jingly
- |
  jingoism
- |
  jingoist
- |
  jingoistic
- |
  Jinnah
- |
  jinnee
- |
  jinni
- |
  jinricksha
- |
  jinrikisha
- |
  jinriksha
- |
  jinxed
- |
  Jinzhou
- |
  jitney
- |
  jitter
- |
  jitterbug
- |
  jitterbugger
- |
  jitteriness
- |
  jitters
- |
  jittery
- |
  jiujitsu
- |
  jiver
- |
  jivey
- |
  Joann
- |
  Joanna
- |
  Joanne
- |
  jobber
- |
  jobholder
- |
  jobless
- |
  joblessness
- |
  Jocasta
- |
  Jocelin
- |
  Jocelyn
- |
  jockey
- |
  jockstrap
- |
  jocose
- |
  jocosely
- |
  jocoseness
- |
  jocosity
- |
  jocular
- |
  jocularity
- |
  jocularly
- |
  jocund
- |
  jocundity
- |
  jocundly
- |
  Jodhpur
- |
  jodhpur
- |
  jodhpurs
- |
  Jodie
- |
  jogger
- |
  jogging
- |
  joggle
- |
  Jogjakarta
- |
  Johanna
- |
  Johannesburg
- |
  johnny
- |
  johnnycake
- |
  Johns
- |
  Johnson
- |
  joinder
- |
  joiner
- |
  joinery
- |
  joint
- |
  jointed
- |
  jointly
- |
  joist
- |
  jojoba
- |
  joker
- |
  jokester
- |
  jokey
- |
  jokingly
- |
  Jolene
- |
  Joliet
- |
  Jolliet
- |
  jollily
- |
  jolliness
- |
  jollity
- |
  jolly
- |
  Jolson
- |
  jolter
- |
  jolty
- |
  Jonah
- |
  Jonas
- |
  Jonathan
- |
  Jones
- |
  jongleur
- |
  jonquil
- |
  Jonson
- |
  Joplin
- |
  Jordan
- |
  Jordanian
- |
  Josef
- |
  Joseph
- |
  Josephine
- |
  Josephus
- |
  josher
- |
  Joshua
- |
  jostle
- |
  jostler
- |
  Josue
- |
  jotter
- |
  jotting
- |
  joule
- |
  jounce
- |
  jouncy
- |
  journal
- |
  journalese
- |
  journalism
- |
  journalist
- |
  journalistic
- |
  journey
- |
  journeyer
- |
  journeyman
- |
  joust
- |
  jouster
- |
  jousting
- |
  jovial
- |
  joviality
- |
  jovially
- |
  jowls
- |
  jowly
- |
  Joyce
- |
  Joycean
- |
  joyful
- |
  joyfully
- |
  joyfulness
- |
  joyless
- |
  joylessly
- |
  joylessness
- |
  joyous
- |
  joyously
- |
  joyousness
- |
  joyridden
- |
  joyride
- |
  joyrider
- |
  joyriding
- |
  joyrode
- |
  joystick
- |
  Juanita
- |
  Juarez
- |
  jubilance
- |
  jubilant
- |
  jubilantly
- |
  jubilation
- |
  jubilee
- |
  Judaea
- |
  Judah
- |
  Judaic
- |
  Judaical
- |
  Judaism
- |
  Judas
- |
  Judea
- |
  Judean
- |
  judge
- |
  judgement
- |
  Judges
- |
  judgeship
- |
  judging
- |
  judgment
- |
  judgmental
- |
  judgmentally
- |
  judicatory
- |
  judicature
- |
  judicial
- |
  judicially
- |
  judiciary
- |
  judicious
- |
  judiciously
- |
  Judie
- |
  Judith
- |
  judoist
- |
  Judson
- |
  Juggernaut
- |
  juggernaut
- |
  juggle
- |
  juggler
- |
  jugglery
- |
  juggling
- |
  Jugoslav
- |
  Jugoslavia
- |
  Jugoslavian
- |
  jugular
- |
  juice
- |
  juiced
- |
  juicer
- |
  juicily
- |
  juiciness
- |
  juicy
- |
  jujitsu
- |
  jujube
- |
  jujutsu
- |
  jukebox
- |
  julep
- |
  Jules
- |
  Julia
- |
  Julian
- |
  Juliana
- |
  Juliann
- |
  Julianne
- |
  Julie
- |
  Julien
- |
  julienne
- |
  Juliet
- |
  Julius
- |
  Julundur
- |
  Jumada
- |
  jumble
- |
  jumbo
- |
  Jumna
- |
  jumper
- |
  jumpers
- |
  jumpily
- |
  jumpiness
- |
  jumps
- |
  jumpsuit
- |
  jumpy
- |
  junco
- |
  junction
- |
  junctional
- |
  juncture
- |
  Juneau
- |
  Jungfrau
- |
  Jungian
- |
  jungle
- |
  junglegym
- |
  jungly
- |
  Junior
- |
  junior
- |
  juniper
- |
  Junker
- |
  junker
- |
  junket
- |
  junketeer
- |
  junketer
- |
  junketing
- |
  junkie
- |
  junky
- |
  junkyard
- |
  junta
- |
  junto
- |
  Jupiter
- |
  Jurassic
- |
  juridic
- |
  juridical
- |
  juridically
- |
  jurisdiction
- |
  jurisprudent
- |
  jurist
- |
  juristic
- |
  juristical
- |
  juror
- |
  jussive
- |
  justice
- |
  justifiable
- |
  justifiably
- |
  justified
- |
  justify
- |
  Justin
- |
  Justina
- |
  Justine
- |
  Justinian
- |
  justly
- |
  justness
- |
  Jutland
- |
  Juvenal
- |
  juvenescence
- |
  juvenescent
- |
  juvenile
- |
  juvenilely
- |
  juvenileness
- |
  juvenilia
- |
  juvenility
- |
  juvenilize
- |
  juvenilized
- |
  juxtapose
- |
  Kaaren
- |
  Kabbala
- |
  Kabbalah
- |
  kabbalah
- |
  Kabbalism
- |
  kabbalism
- |
  Kabbalist
- |
  kabbalist
- |
  Kabbalistic
- |
  kabbalistic
- |
  kabob
- |
  Kabuki
- |
  kabuki
- |
  Kabul
- |
  kachina
- |
  Kadar
- |
  Kaddish
- |
  kaddish
- |
  kaffeeklatch
- |
  Kaffir
- |
  kaffiyeh
- |
  kafir
- |
  Kafka
- |
  Kafkaesque
- |
  kaftan
- |
  Kagoshima
- |
  kahuna
- |
  Kaiser
- |
  kaiser
- |
  Kaiserin
- |
  kaisership
- |
  Kalahari
- |
  Kalamazoo
- |
  kaleidoscope
- |
  kalends
- |
  Kalgan
- |
  Kalimantan
- |
  kalimba
- |
  Kalinin
- |
  Kaliningrad
- |
  Kaluga
- |
  Kalyan
- |
  kamaaina
- |
  Kamchatka
- |
  Kamehameha
- |
  Kamet
- |
  kamikaze
- |
  Kampala
- |
  Kampuchea
- |
  Kampuchean
- |
  kanaka
- |
  Kananga
- |
  Kanchenjunga
- |
  Kandinski
- |
  Kandinsky
- |
  kangaroo
- |
  Kanpur
- |
  Kansan
- |
  Kansas
- |
  Kantian
- |
  Kaohsiung
- |
  kaolin
- |
  kaoline
- |
  kapok
- |
  kappa
- |
  kaput
- |
  kaputt
- |
  Karachi
- |
  Karaganda
- |
  Karaj
- |
  karakul
- |
  karaoke
- |
  karat
- |
  karate
- |
  Karelia
- |
  Karelian
- |
  Karen
- |
  Karin
- |
  Karla
- |
  Karlsruhe
- |
  karma
- |
  karmic
- |
  karmically
- |
  Karol
- |
  Karolyn
- |
  Karoo
- |
  Karroo
- |
  karst
- |
  karstic
- |
  karstify
- |
  karyotype
- |
  Kashmir
- |
  Kashmiri
- |
  katabatic
- |
  katakana
- |
  Katharine
- |
  Katherine
- |
  Kathiawar
- |
  Kathleen
- |
  Kathmandu
- |
  Kathryn
- |
  Kathy
- |
  Katie
- |
  Katmandu
- |
  Katowice
- |
  Kattegat
- |
  katydid
- |
  Kauai
- |
  Kaunas
- |
  Kaunda
- |
  Kawabata
- |
  Kawasaki
- |
  kayak
- |
  kayaker
- |
  Kayseri
- |
  Kazakh
- |
  Kazakhstan
- |
  Kazan
- |
  kazoo
- |
  Keats
- |
  Keatsian
- |
  kebab
- |
  kebob
- |
  kedge
- |
  keelboat
- |
  keeled
- |
  keelhaul
- |
  Keelung
- |
  keener
- |
  keenly
- |
  keenness
- |
  keeper
- |
  keeping
- |
  keepsake
- |
  Keewatin
- |
  keffiyeh
- |
  kegler
- |
  Keith
- |
  Keller
- |
  Kellogg
- |
  Kelly
- |
  Kelvin
- |
  kelvin
- |
  Kemerovo
- |
  Kempis
- |
  Kenai
- |
  Kendall
- |
  Kennedy
- |
  kennel
- |
  kennels
- |
  Kenneth
- |
  Kenny
- |
  kente
- |
  Kentish
- |
  Kenton
- |
  Kentuckian
- |
  Kentucky
- |
  Kenya
- |
  Kenyan
- |
  Kenyatta
- |
  Keokuk
- |
  Kepler
- |
  keratin
- |
  keratinous
- |
  kerchief
- |
  kerchieves
- |
  Kerensky
- |
  Kerman
- |
  kermes
- |
  kermis
- |
  Kermit
- |
  kerne
- |
  kernel
- |
  kerning
- |
  kerosene
- |
  kerosine
- |
  Kerouac
- |
  Kerry
- |
  kestrel
- |
  ketch
- |
  ketchup
- |
  ketone
- |
  kettle
- |
  kettledrum
- |
  Kevin
- |
  Kevlar
- |
  keyboard
- |
  keyboarder
- |
  keyboardist
- |
  keycard
- |
  keyhole
- |
  Keynes
- |
  Keynesian
- |
  Keynesianism
- |
  keynote
- |
  keynoter
- |
  keypad
- |
  keypunch
- |
  keypuncher
- |
  keystone
- |
  keystroke
- |
  keyword
- |
  Khabarovsk
- |
  Khachaturian
- |
  khaki
- |
  khakis
- |
  Khalid
- |
  khanate
- |
  Kharkiv
- |
  Kharkov
- |
  Khartoum
- |
  Khayyam
- |
  khedive
- |
  Kherson
- |
  Khmer
- |
  Khoisan
- |
  Khomeini
- |
  khoum
- |
  Khrushchev
- |
  Khufu
- |
  Khulna
- |
  Khyber
- |
  kibble
- |
  kibbutz
- |
  kibbutzim
- |
  kibitz
- |
  kibitzer
- |
  kibosh
- |
  Kickapoo
- |
  kickback
- |
  kicker
- |
  kickoff
- |
  kicks
- |
  kickshaw
- |
  kickstand
- |
  kickstart
- |
  kicky
- |
  kidder
- |
  kiddie
- |
  kiddingly
- |
  kiddish
- |
  kiddo
- |
  kiddy
- |
  kidnap
- |
  kidnaper
- |
  kidnapper
- |
  kidnapping
- |
  kidney
- |
  kidskin
- |
  kielbasa
- |
  kielbasi
- |
  kielbasy
- |
  Kierkegaard
- |
  Kievan
- |
  Kigali
- |
  Kikuyu
- |
  Kilauea
- |
  Kilimanjaro
- |
  killdeer
- |
  killer
- |
  killing
- |
  killjoy
- |
  kilobit
- |
  kilobyte
- |
  kilocalorie
- |
  kilocycle
- |
  kilogram
- |
  kilogramme
- |
  kilohertz
- |
  kiloliter
- |
  kilometer
- |
  kilometre
- |
  kilometric
- |
  kiloton
- |
  kilovolt
- |
  kilowatt
- |
  kilter
- |
  Kimberly
- |
  kimchi
- |
  kimono
- |
  kinaesthesia
- |
  kinda
- |
  kindergarten
- |
  kindhearted
- |
  kindle
- |
  kindliness
- |
  kindling
- |
  kindly
- |
  kindness
- |
  kindred
- |
  kinema
- |
  kinematic
- |
  kinematical
- |
  kinematics
- |
  kinescope
- |
  kinesics
- |
  kinesiology
- |
  kinesthesia
- |
  kinesthetic
- |
  kinetic
- |
  kinetically
- |
  kinetics
- |
  kinfolk
- |
  kinfolks
- |
  kingbolt
- |
  kingdom
- |
  kingfisher
- |
  kingless
- |
  kingliness
- |
  kingly
- |
  kingpin
- |
  Kings
- |
  kingship
- |
  Kingston
- |
  Kingstown
- |
  kinkajou
- |
  kinkily
- |
  kinkiness
- |
  kinky
- |
  Kinsey
- |
  kinsfolk
- |
  Kinshasa
- |
  kinship
- |
  kinsman
- |
  kinswoman
- |
  kiosk
- |
  Kiowa
- |
  Kipling
- |
  kipper
- |
  Kirby
- |
  Kirghiz
- |
  Kirghizia
- |
  Kiribati
- |
  kirigami
- |
  Kirin
- |
  Kirkuk
- |
  Kirkwall
- |
  Kirov
- |
  kirsch
- |
  kirtle
- |
  Kisangani
- |
  Kishinev
- |
  Kishinyov
- |
  Kislev
- |
  kismet
- |
  kissable
- |
  kisser
- |
  Kissinger
- |
  Kitakyushu
- |
  kitbag
- |
  kitchen
- |
  Kitchener
- |
  kitchenet
- |
  kitchenette
- |
  kitchenware
- |
  kitsch
- |
  kitschiness
- |
  kitschy
- |
  kitten
- |
  kittenish
- |
  kittenishly
- |
  Kitty
- |
  kitty
- |
  kittycat
- |
  Kitwe
- |
  kiwifruit
- |
  Klamath
- |
  klatch
- |
  klatsch
- |
  Klaus
- |
  Kleenex
- |
  kleptomania
- |
  kleptomaniac
- |
  Klondike
- |
  klutz
- |
  klutziness
- |
  klutzy
- |
  knack
- |
  knackwurst
- |
  knapsack
- |
  knave
- |
  knavery
- |
  knavish
- |
  knavishly
- |
  knavishness
- |
  knead
- |
  kneader
- |
  kneading
- |
  kneecap
- |
  kneed
- |
  kneehole
- |
  kneel
- |
  knell
- |
  knelt
- |
  Knesset
- |
  knickers
- |
  knickknack
- |
  knife
- |
  knight
- |
  knighthood
- |
  knightly
- |
  knish
- |
  knitter
- |
  knitting
- |
  knitwear
- |
  knives
- |
  knobbed
- |
  knobby
- |
  knoblike
- |
  knock
- |
  knockdown
- |
  knocker
- |
  knocking
- |
  knockoff
- |
  knockout
- |
  knockwurst
- |
  knoll
- |
  Knossus
- |
  knothole
- |
  knottiness
- |
  knotty
- |
  knout
- |
  knowable
- |
  knower
- |
  knowhow
- |
  knowing
- |
  knowingly
- |
  knowledge
- |
  known
- |
  Knoxville
- |
  knuckle
- |
  knucklebone
- |
  knucklehead
- |
  knurl
- |
  knurled
- |
  knurly
- |
  koala
- |
  Koblenz
- |
  Kodaly
- |
  Kodiak
- |
  Koestler
- |
  kohlrabi
- |
  kolinsky
- |
  Kolwesi
- |
  Kolyma
- |
  Komsomolsk
- |
  Konya
- |
  kookaburra
- |
  kookie
- |
  kookiness
- |
  kooky
- |
  kopeck
- |
  kopek
- |
  Koran
- |
  Koranic
- |
  Korea
- |
  Korean
- |
  koruna
- |
  Kosciusko
- |
  Kosciuszko
- |
  kosher
- |
  Kosice
- |
  Kosovar
- |
  Kosovo
- |
  Kossuth
- |
  Kosygin
- |
  Kotah
- |
  Kowloon
- |
  kowtow
- |
  kowtower
- |
  kraal
- |
  Krakatau
- |
  Krakatoa
- |
  Krakow
- |
  Krasnodar
- |
  Krasnoyarsk
- |
  kraut
- |
  Kremlin
- |
  kremlin
- |
  Kremlinology
- |
  krill
- |
  Krishna
- |
  Kristin
- |
  Kristine
- |
  krona
- |
  krone
- |
  kroner
- |
  kronor
- |
  kronur
- |
  kroon
- |
  krooni
- |
  Krugerrand
- |
  krugerrand
- |
  krypton
- |
  Kubrick
- |
  kuchen
- |
  kudos
- |
  kudzu
- |
  Kueiyang
- |
  Kuibyshev
- |
  kulak
- |
  Kumamoto
- |
  Kumasi
- |
  kummel
- |
  kumquat
- |
  Kunlun
- |
  Kunming
- |
  Kuomintang
- |
  Kurdish
- |
  Kurdistan
- |
  Kuril
- |
  Kurile
- |
  Kurilian
- |
  Kurosawa
- |
  Kursk
- |
  kurus
- |
  Kuwait
- |
  Kuwaiti
- |
  Kuybyshev
- |
  Kuzbas
- |
  Kuzbass
- |
  kvetch
- |
  kvetcher
- |
  kwacha
- |
  Kwajalein
- |
  Kwakiutl
- |
  Kwangchow
- |
  Kwangju
- |
  Kwanza
- |
  kwanza
- |
  Kwanzaa
- |
  kwashiorkor
- |
  Kweiyang
- |
  Kyoto
- |
  Kyrgyz
- |
  Kyrgyzstan
- |
  Kyushu
- |
  label
- |
  labeler
- |
  labeller
- |
  labia
- |
  labial
- |
  labialize
- |
  labially
- |
  labile
- |
  lability
- |
  labium
- |
  labor
- |
  laboratory
- |
  labored
- |
  laborer
- |
  laborious
- |
  laboriously
- |
  laborsaving
- |
  labour
- |
  labourer
- |
  Labrador
- |
  Labradorean
- |
  Labradorian
- |
  labradorite
- |
  labret
- |
  laburnum
- |
  Labyrinth
- |
  labyrinth
- |
  labyrinthian
- |
  labyrinthine
- |
  Laccadive
- |
  Lacedaemon
- |
  lacer
- |
  lacerate
- |
  lacerated
- |
  laceration
- |
  Lacerta
- |
  laces
- |
  lacewing
- |
  lacework
- |
  Lachesis
- |
  lachrymal
- |
  lachrymose
- |
  lachrymosely
- |
  lachrymosity
- |
  laciness
- |
  lackey
- |
  lacking
- |
  lackluster
- |
  lacklustre
- |
  Laconia
- |
  Laconian
- |
  laconic
- |
  laconically
- |
  laconicism
- |
  laconism
- |
  lacquer
- |
  lacquered
- |
  lacquey
- |
  lacrimal
- |
  lacrimation
- |
  lacrosse
- |
  lacrymal
- |
  lactate
- |
  lactation
- |
  lactational
- |
  lacteal
- |
  lactic
- |
  lactose
- |
  lacuna
- |
  lacunae
- |
  lacunal
- |
  lacunary
- |
  lacunate
- |
  lacunose
- |
  lacustrine
- |
  ladder
- |
  laddie
- |
  laden
- |
  lading
- |
  Ladino
- |
  ladle
- |
  ladler
- |
  Ladoga
- |
  ladybird
- |
  ladybug
- |
  ladyfinger
- |
  ladylike
- |
  ladylove
- |
  Ladyship
- |
  ladyship
- |
  laetrile
- |
  Lafayette
- |
  Lafitte
- |
  LaFollette
- |
  lager
- |
  laggard
- |
  laggardly
- |
  laggardness
- |
  lagger
- |
  lagging
- |
  lagnappe
- |
  lagniappe
- |
  lagoon
- |
  lagoonal
- |
  Lagos
- |
  Lahore
- |
  laical
- |
  laically
- |
  laird
- |
  lairdship
- |
  laity
- |
  Laius
- |
  Lakehurst
- |
  Lakewood
- |
  Lakota
- |
  lalapalooza
- |
  lallygag
- |
  Lamaism
- |
  Lamaist
- |
  Lamaistic
- |
  Lamar
- |
  Lamarck
- |
  lamasery
- |
  Lamaze
- |
  lambada
- |
  lambast
- |
  lambaste
- |
  lambda
- |
  lambency
- |
  lambent
- |
  lambently
- |
  Lambeth
- |
  lambkin
- |
  lambskin
- |
  lamebrain
- |
  lamella
- |
  lamellae
- |
  lamellar
- |
  lamellate
- |
  lamely
- |
  lameness
- |
  lament
- |
  lamentable
- |
  lamentably
- |
  lamentation
- |
  Lamentations
- |
  lamenter
- |
  lamia
- |
  lamina
- |
  laminable
- |
  laminae
- |
  laminal
- |
  laminar
- |
  laminate
- |
  laminated
- |
  lamination
- |
  laminator
- |
  laminose
- |
  lampblack
- |
  lamplighter
- |
  lampoon
- |
  lampooner
- |
  lampoonist
- |
  lamppost
- |
  lamprey
- |
  lampshade
- |
  Lanai
- |
  lanai
- |
  Lancashire
- |
  Lancaster
- |
  Lancastrian
- |
  Lance
- |
  lance
- |
  Lancelot
- |
  lancer
- |
  lancet
- |
  lanceted
- |
  Lanchou
- |
  Lanchow
- |
  landau
- |
  landed
- |
  lander
- |
  landfall
- |
  landfill
- |
  landform
- |
  landholder
- |
  landholding
- |
  landing
- |
  landlady
- |
  landless
- |
  landlocked
- |
  landlord
- |
  landlubber
- |
  landlubberly
- |
  landmark
- |
  landmass
- |
  landowner
- |
  landowning
- |
  landscape
- |
  landscaper
- |
  landscaping
- |
  landslide
- |
  landsman
- |
  landward
- |
  landwards
- |
  Langland
- |
  Langley
- |
  language
- |
  Languedoc
- |
  languid
- |
  languidly
- |
  languidness
- |
  languish
- |
  languisher
- |
  languor
- |
  languorous
- |
  languorously
- |
  laniard
- |
  lankily
- |
  lankiness
- |
  lankly
- |
  lankness
- |
  lanky
- |
  Lanny
- |
  lanolin
- |
  Lansing
- |
  lantana
- |
  lantern
- |
  lanthanide
- |
  lanthanum
- |
  lanyard
- |
  Lanzhou
- |
  Laocoon
- |
  Laodicean
- |
  Laotian
- |
  Laozi
- |
  laparoscope
- |
  laparoscopic
- |
  laparoscopy
- |
  lapboard
- |
  lapdog
- |
  lapel
- |
  lapeled
- |
  lapelled
- |
  lapful
- |
  lapidary
- |
  lapin
- |
  Laplace
- |
  Lapland
- |
  Laplander
- |
  lappet
- |
  lapping
- |
  Lappish
- |
  lapse
- |
  lapser
- |
  laptop
- |
  lapwing
- |
  larboard
- |
  larcenist
- |
  larcenous
- |
  larceny
- |
  larch
- |
  larder
- |
  lardy
- |
  Laredo
- |
  lares
- |
  large
- |
  largehearted
- |
  largely
- |
  largeness
- |
  largess
- |
  largesse
- |
  largish
- |
  Largo
- |
  largo
- |
  lariat
- |
  larker
- |
  larkish
- |
  larkspur
- |
  Larne
- |
  Larousse
- |
  Larry
- |
  larva
- |
  larvae
- |
  larval
- |
  larvicide
- |
  laryngeal
- |
  larynges
- |
  laryngitic
- |
  laryngitis
- |
  larynx
- |
  lasagna
- |
  lasagne
- |
  lascar
- |
  lascivious
- |
  lasciviously
- |
  laser
- |
  lasher
- |
  lashings
- |
  lassie
- |
  lassitude
- |
  lasso
- |
  lassoer
- |
  lasting
- |
  lastingly
- |
  lastingness
- |
  lastly
- |
  Latakia
- |
  latch
- |
  latchet
- |
  latchkey
- |
  latchstring
- |
  latecomer
- |
  lateen
- |
  lately
- |
  latency
- |
  lateness
- |
  latent
- |
  latently
- |
  later
- |
  lateral
- |
  laterally
- |
  latest
- |
  latex
- |
  lathe
- |
  lather
- |
  latherer
- |
  lathery
- |
  latices
- |
  Latin
- |
  Latina
- |
  Latino
- |
  latino
- |
  latish
- |
  latitude
- |
  latitudes
- |
  latitudinal
- |
  Latium
- |
  latke
- |
  latrine
- |
  latte
- |
  latter
- |
  latterly
- |
  lattice
- |
  latticed
- |
  latticework
- |
  Latvia
- |
  Latvian
- |
  laudability
- |
  laudable
- |
  laudableness
- |
  laudably
- |
  laudanum
- |
  laudation
- |
  laudatory
- |
  lauded
- |
  lauder
- |
  laugh
- |
  laughable
- |
  laughably
- |
  laugher
- |
  laughing
- |
  laughingly
- |
  laughs
- |
  laughter
- |
  launch
- |
  launcher
- |
  launchpad
- |
  launder
- |
  launderer
- |
  launderette
- |
  laundress
- |
  Laundromat
- |
  laundromat
- |
  laundry
- |
  laundryman
- |
  laundrywoman
- |
  Laura
- |
  laureate
- |
  laureateship
- |
  Laurel
- |
  laurel
- |
  laurels
- |
  Lauren
- |
  Laurence
- |
  Laurentian
- |
  Laurie
- |
  Lausanne
- |
  lavage
- |
  Laval
- |
  lavalier
- |
  lavaliere
- |
  lavash
- |
  lavatory
- |
  lavender
- |
  Lavern
- |
  Laverne
- |
  Lavinia
- |
  lavish
- |
  lavisher
- |
  lavishly
- |
  lavishness
- |
  Lavoisier
- |
  lawbreaker
- |
  lawbreaking
- |
  lawful
- |
  lawfully
- |
  lawfulness
- |
  lawgiver
- |
  lawless
- |
  lawlessly
- |
  lawlessness
- |
  lawmaker
- |
  lawmaking
- |
  lawman
- |
  lawnmower
- |
  Lawrence
- |
  lawrencium
- |
  lawsuit
- |
  lawyer
- |
  lawyerly
- |
  laxation
- |
  laxative
- |
  laxity
- |
  laxly
- |
  laxness
- |
  Layamon
- |
  layaway
- |
  layer
- |
  layered
- |
  layette
- |
  layman
- |
  layoff
- |
  layout
- |
  layover
- |
  laypeople
- |
  layperson
- |
  Layton
- |
  laywoman
- |
  lazar
- |
  Lazarus
- |
  lazily
- |
  laziness
- |
  lazybones
- |
  leach
- |
  leacher
- |
  leaded
- |
  leaden
- |
  leadenly
- |
  leadenness
- |
  leader
- |
  leaderless
- |
  leadership
- |
  leading
- |
  leafage
- |
  leafed
- |
  leafhopper
- |
  leafiness
- |
  leafless
- |
  leaflet
- |
  leafstalk
- |
  leafy
- |
  league
- |
  leakage
- |
  leaker
- |
  Leakey
- |
  leakiness
- |
  leaky
- |
  Leander
- |
  leaner
- |
  leaning
- |
  leanly
- |
  Leanne
- |
  leanness
- |
  leant
- |
  leaper
- |
  leapfrog
- |
  leapt
- |
  learn
- |
  learned
- |
  learnedly
- |
  learnedness
- |
  learner
- |
  learning
- |
  learnt
- |
  Leary
- |
  lease
- |
  leaseback
- |
  leasehold
- |
  leaseholder
- |
  leaser
- |
  leash
- |
  least
- |
  leastways
- |
  leastwise
- |
  leather
- |
  leatherback
- |
  leatherette
- |
  leatheriness
- |
  leathern
- |
  leatherneck
- |
  leathery
- |
  leave
- |
  leaved
- |
  leaven
- |
  leavening
- |
  leaver
- |
  leaves
- |
  leavings
- |
  Lebanese
- |
  Lebanon
- |
  lecher
- |
  lecherous
- |
  lecherously
- |
  lechery
- |
  lecithin
- |
  lectern
- |
  lection
- |
  lectionary
- |
  lector
- |
  lecture
- |
  lecturer
- |
  lectureship
- |
  lederhosen
- |
  ledge
- |
  ledger
- |
  leech
- |
  Leeds
- |
  leerily
- |
  leeriness
- |
  leeringly
- |
  leery
- |
  Leeuwenhoek
- |
  leeward
- |
  leeway
- |
  Leftism
- |
  leftism
- |
  leftist
- |
  leftmost
- |
  leftover
- |
  leftovers
- |
  lefty
- |
  legacy
- |
  legal
- |
  legalese
- |
  legalise
- |
  legalism
- |
  legalist
- |
  legalistic
- |
  legality
- |
  legalization
- |
  legalize
- |
  legally
- |
  legate
- |
  legatee
- |
  legateship
- |
  legatine
- |
  legation
- |
  legationary
- |
  legato
- |
  legend
- |
  legendarily
- |
  legendary
- |
  legerdemain
- |
  legged
- |
  leggin
- |
  legginess
- |
  legging
- |
  leggings
- |
  leggy
- |
  Leghorn
- |
  leghorn
- |
  legibility
- |
  legible
- |
  legibleness
- |
  legibly
- |
  legion
- |
  legionary
- |
  legionnaire
- |
  legions
- |
  legislate
- |
  legislation
- |
  legislative
- |
  legislator
- |
  legislature
- |
  legit
- |
  legitimacy
- |
  legitimate
- |
  legitimately
- |
  legitimation
- |
  legitimatize
- |
  legitimise
- |
  legitimism
- |
  legitimist
- |
  legitimize
- |
  legless
- |
  legman
- |
  Legree
- |
  legroom
- |
  legume
- |
  leguminous
- |
  legwork
- |
  Leibnitz
- |
  Leibniz
- |
  Leicester
- |
  Leiden
- |
  Leigh
- |
  Leighton
- |
  Leila
- |
  Leinster
- |
  Leipzig
- |
  leisure
- |
  leisured
- |
  leisurely
- |
  leisurewear
- |
  leitmotif
- |
  leitmotiv
- |
  Leland
- |
  Lelia
- |
  Leman
- |
  lemma
- |
  lemmata
- |
  lemming
- |
  Lemnos
- |
  lemon
- |
  lemonade
- |
  lemony
- |
  lempira
- |
  Lemuel
- |
  lemur
- |
  lender
- |
  lending
- |
  length
- |
  lengthen
- |
  lengthily
- |
  lengthiness
- |
  lengths
- |
  lengthways
- |
  lengthwise
- |
  lengthy
- |
  lenience
- |
  leniency
- |
  lenient
- |
  leniently
- |
  Lenin
- |
  Leningrad
- |
  Leninism
- |
  Leninist
- |
  lenitive
- |
  lenity
- |
  Lennon
- |
  Lenora
- |
  Lenore
- |
  Lenten
- |
  lenten
- |
  lentil
- |
  lento
- |
  Leona
- |
  Leonard
- |
  Leoncavallo
- |
  leone
- |
  leonine
- |
  Leonora
- |
  Leonore
- |
  leopard
- |
  Leopold
- |
  leotard
- |
  leotarded
- |
  leotards
- |
  leper
- |
  lepidoptery
- |
  leprechaun
- |
  leprosy
- |
  leprous
- |
  leptin
- |
  lepton
- |
  leptonic
- |
  Lepus
- |
  Lerner
- |
  Leroy
- |
  Lerwick
- |
  lesbian
- |
  lesbianism
- |
  lesion
- |
  Lesley
- |
  Leslie
- |
  Lesotho
- |
  lessee
- |
  lesseeship
- |
  lessen
- |
  lessening
- |
  Lesseps
- |
  lesser
- |
  Lessing
- |
  lesson
- |
  lessor
- |
  Lester
- |
  letdown
- |
  lethal
- |
  lethality
- |
  lethally
- |
  lethargic
- |
  lethargy
- |
  Lethe
- |
  lethe
- |
  Letitia
- |
  letter
- |
  lettered
- |
  letterer
- |
  letterhead
- |
  lettering
- |
  letterpress
- |
  letters
- |
  Lettish
- |
  lettuce
- |
  letup
- |
  leucocyte
- |
  leukaemia
- |
  leukemia
- |
  leukemic
- |
  leukocyte
- |
  leukocytic
- |
  Levant
- |
  Levantine
- |
  levee
- |
  level
- |
  leveler
- |
  levelheaded
- |
  leveller
- |
  levelly
- |
  levelness
- |
  lever
- |
  leverage
- |
  leveraged
- |
  leviable
- |
  Leviathan
- |
  leviathan
- |
  levier
- |
  levies
- |
  Levis
- |
  levis
- |
  levitate
- |
  levitation
- |
  levitator
- |
  Leviticus
- |
  Levittown
- |
  levity
- |
  lewdly
- |
  lewdness
- |
  Lewes
- |
  Lewis
- |
  Lewisham
- |
  Lewiston
- |
  lexica
- |
  lexical
- |
  lexically
- |
  lexicography
- |
  lexicon
- |
  Lexington
- |
  lexis
- |
  Leyden
- |
  Leyte
- |
  Lhasa
- |
  liabilities
- |
  liability
- |
  liable
- |
  liaise
- |
  liaison
- |
  liana
- |
  libation
- |
  Libby
- |
  libel
- |
  libeler
- |
  libelist
- |
  libeller
- |
  libellous
- |
  libelous
- |
  libelously
- |
  Liberal
- |
  liberal
- |
  liberalise
- |
  liberalism
- |
  liberalist
- |
  liberalistic
- |
  liberality
- |
  liberalize
- |
  liberally
- |
  liberalness
- |
  liberate
- |
  liberated
- |
  liberation
- |
  liberator
- |
  Liberia
- |
  Liberian
- |
  libertarian
- |
  liberties
- |
  libertinage
- |
  libertine
- |
  libertinism
- |
  Liberty
- |
  liberty
- |
  libidinal
- |
  libidinally
- |
  libidinous
- |
  libidinously
- |
  libido
- |
  Libra
- |
  librarian
- |
  library
- |
  libretti
- |
  librettist
- |
  libretto
- |
  Libreville
- |
  Libya
- |
  Libyan
- |
  licence
- |
  licensable
- |
  license
- |
  licensed
- |
  licensee
- |
  licenser
- |
  licensing
- |
  licente
- |
  licentiate
- |
  licentious
- |
  licentiously
- |
  lichee
- |
  lichen
- |
  lichened
- |
  lichenology
- |
  lichenous
- |
  Lichtenstein
- |
  licit
- |
  licitly
- |
  licitness
- |
  licker
- |
  licking
- |
  lickspittle
- |
  licorice
- |
  lidded
- |
  lidocaine
- |
  lieder
- |
  Liege
- |
  liege
- |
  lieutenancy
- |
  Lieutenant
- |
  lieutenant
- |
  lifebelt
- |
  lifeblood
- |
  lifeboat
- |
  lifebuoy
- |
  lifecare
- |
  lifeguard
- |
  lifeless
- |
  lifelessly
- |
  lifelessness
- |
  lifelike
- |
  lifeline
- |
  lifelong
- |
  lifer
- |
  Lifesaver
- |
  lifesaver
- |
  lifesaving
- |
  lifestyle
- |
  lifetime
- |
  lifework
- |
  Liffey
- |
  liftable
- |
  lifter
- |
  liftoff
- |
  ligament
- |
  ligate
- |
  ligation
- |
  ligature
- |
  light
- |
  lighted
- |
  lighten
- |
  lightener
- |
  lighter
- |
  lightface
- |
  lightfaced
- |
  lightheaded
- |
  lighthearted
- |
  lighthouse
- |
  lighting
- |
  lightish
- |
  lightly
- |
  lightness
- |
  lightning
- |
  lightproof
- |
  lights
- |
  lightship
- |
  lightsome
- |
  lightweight
- |
  lightyear
- |
  ligneous
- |
  lignin
- |
  lignite
- |
  lignitic
- |
  ligroin
- |
  Liguria
- |
  Ligurian
- |
  likability
- |
  likable
- |
  likableness
- |
  likably
- |
  likeability
- |
  likeable
- |
  likeableness
- |
  likeably
- |
  likelihood
- |
  likely
- |
  liken
- |
  likeness
- |
  likes
- |
  likewise
- |
  liking
- |
  likuta
- |
  lilac
- |
  lilangeni
- |
  Liliuokalani
- |
  Lille
- |
  Lillian
- |
  Lillie
- |
  Lilliput
- |
  Lilliputian
- |
  lilliputian
- |
  Lilongwe
- |
  lilting
- |
  Limavady
- |
  limber
- |
  limberness
- |
  limbic
- |
  limbless
- |
  Limbo
- |
  limbo
- |
  Limburger
- |
  limeade
- |
  limelight
- |
  limerick
- |
  limestone
- |
  Limey
- |
  limit
- |
  limitable
- |
  limitation
- |
  limited
- |
  limitedly
- |
  limiter
- |
  limiting
- |
  limitless
- |
  limits
- |
  limner
- |
  limnology
- |
  Limoges
- |
  limonite
- |
  limonitic
- |
  limousine
- |
  limpet
- |
  limpid
- |
  limpidity
- |
  limpidly
- |
  limpidness
- |
  limply
- |
  limpness
- |
  Limpopo
- |
  linage
- |
  linchpin
- |
  Lincoln
- |
  Lincolnshire
- |
  Linda
- |
  Lindbergh
- |
  linden
- |
  Lindsay
- |
  Lindsey
- |
  lineage
- |
  lineal
- |
  lineally
- |
  lineament
- |
  lineaments
- |
  linear
- |
  linearity
- |
  linearly
- |
  lineation
- |
  linebacker
- |
  lined
- |
  lineman
- |
  linen
- |
  linens
- |
  liner
- |
  linerless
- |
  lines
- |
  linesman
- |
  lineup
- |
  linger
- |
  lingerer
- |
  lingerie
- |
  lingering
- |
  lingeringly
- |
  lingo
- |
  lingual
- |
  lingually
- |
  linguine
- |
  linguini
- |
  linguist
- |
  linguistic
- |
  linguistics
- |
  liniment
- |
  lining
- |
  linkage
- |
  linker
- |
  links
- |
  linkup
- |
  Linnaean
- |
  Linnaeus
- |
  Linnean
- |
  linnet
- |
  linoleum
- |
  linseed
- |
  lintel
- |
  linteled
- |
  lintelled
- |
  linty
- |
  Lionel
- |
  lioness
- |
  lionhearted
- |
  lionization
- |
  lionize
- |
  lionizer
- |
  Lipetsk
- |
  lipid
- |
  lipide
- |
  lipidic
- |
  lipoprotein
- |
  liposuction
- |
  lipotropic
- |
  lipotropin
- |
  lipped
- |
  Lippi
- |
  lippiness
- |
  Lippmann
- |
  lippy
- |
  lipread
- |
  lipreader
- |
  lipreading
- |
  lipstick
- |
  lipsticked
- |
  lipsynch
- |
  liquefaction
- |
  liquefactive
- |
  liquefiable
- |
  liquefier
- |
  liquefy
- |
  liqueur
- |
  liquid
- |
  liquidate
- |
  liquidation
- |
  liquidator
- |
  liquidity
- |
  liquidize
- |
  liquidizer
- |
  liquidness
- |
  liquify
- |
  liquor
- |
  liquorice
- |
  Lisbon
- |
  Lisburn
- |
  lisente
- |
  lisle
- |
  lisper
- |
  lissom
- |
  lissome
- |
  lissomely
- |
  lissomeness
- |
  listee
- |
  listen
- |
  listener
- |
  listenership
- |
  Lister
- |
  listing
- |
  listless
- |
  listlessly
- |
  listlessness
- |
  lists
- |
  listserver
- |
  Liszt
- |
  litany
- |
  litas
- |
  litchi
- |
  liter
- |
  literacy
- |
  literal
- |
  literalism
- |
  literalist
- |
  literalistic
- |
  literality
- |
  literalize
- |
  literally
- |
  literalness
- |
  literarily
- |
  literariness
- |
  literary
- |
  literate
- |
  literately
- |
  literati
- |
  literature
- |
  lithe
- |
  lithely
- |
  litheness
- |
  lithesome
- |
  lithium
- |
  lithograph
- |
  lithographer
- |
  lithographic
- |
  lithography
- |
  lithologic
- |
  lithological
- |
  lithology
- |
  lithosphere
- |
  Lithuania
- |
  Lithuanian
- |
  litigant
- |
  litigate
- |
  litigation
- |
  litigative
- |
  litigator
- |
  litigious
- |
  litigiously
- |
  litmus
- |
  litotes
- |
  litre
- |
  litter
- |
  litterbug
- |
  littered
- |
  litterer
- |
  little
- |
  littleneck
- |
  littleness
- |
  littoral
- |
  liturgical
- |
  liturgically
- |
  liturgist
- |
  Liturgy
- |
  liturgy
- |
  livability
- |
  livable
- |
  livableness
- |
  liveable
- |
  livebearer
- |
  lived
- |
  livelihood
- |
  livelily
- |
  liveliness
- |
  livelong
- |
  lively
- |
  liven
- |
  liver
- |
  liveried
- |
  liverish
- |
  liverishness
- |
  Liverpool
- |
  Liverpudlian
- |
  liverwort
- |
  liverwurst
- |
  livery
- |
  liveryman
- |
  lives
- |
  livestock
- |
  livid
- |
  lividity
- |
  lividly
- |
  lividness
- |
  living
- |
  Livingstone
- |
  Livonia
- |
  Livonian
- |
  Livorno
- |
  livre
- |
  lizard
- |
  Ljubljana
- |
  llama
- |
  llano
- |
  Llewellyn
- |
  Llewelyn
- |
  Lloyd
- |
  loaded
- |
  loader
- |
  loading
- |
  loads
- |
  loadstar
- |
  loadstone
- |
  Loafer
- |
  loafer
- |
  loamy
- |
  loaner
- |
  loansharking
- |
  loanword
- |
  loath
- |
  loathe
- |
  loather
- |
  loathing
- |
  loathingly
- |
  loathsome
- |
  loaves
- |
  lobar
- |
  lobate
- |
  lobber
- |
  lobby
- |
  lobbyer
- |
  lobbying
- |
  lobbyist
- |
  lobed
- |
  lobotomize
- |
  lobotomy
- |
  lobster
- |
  local
- |
  locale
- |
  localised
- |
  locality
- |
  localization
- |
  localize
- |
  localized
- |
  locally
- |
  locate
- |
  located
- |
  locater
- |
  location
- |
  locational
- |
  locative
- |
  locator
- |
  lockable
- |
  lockbox
- |
  Locke
- |
  locked
- |
  locker
- |
  locket
- |
  lockjaw
- |
  locknut
- |
  lockout
- |
  locks
- |
  locksmith
- |
  lockstep
- |
  lockup
- |
  locomotion
- |
  locomotive
- |
  locomotor
- |
  locoweed
- |
  locus
- |
  locust
- |
  locution
- |
  locutionary
- |
  loden
- |
  lodestar
- |
  lodestone
- |
  lodge
- |
  lodgement
- |
  lodger
- |
  lodging
- |
  lodgings
- |
  lodgment
- |
  loess
- |
  Loewe
- |
  Lofoten
- |
  loftily
- |
  loftiness
- |
  lofty
- |
  Logan
- |
  loganberry
- |
  logarithm
- |
  logarithmic
- |
  logbook
- |
  logger
- |
  loggerhead
- |
  loggerheads
- |
  loggia
- |
  logging
- |
  loggy
- |
  logic
- |
  logical
- |
  logicality
- |
  logically
- |
  logicalness
- |
  logician
- |
  login
- |
  loginess
- |
  logistic
- |
  logistical
- |
  logistically
- |
  logistics
- |
  logjam
- |
  logon
- |
  logotype
- |
  logroller
- |
  logrolling
- |
  loincloth
- |
  loins
- |
  Loire
- |
  loiter
- |
  loiterer
- |
  loitering
- |
  lollapaloosa
- |
  lollapalooza
- |
  loller
- |
  lollipop
- |
  lollygag
- |
  lollypop
- |
  Lombard
- |
  Lombardy
- |
  London
- |
  Londonderry
- |
  Londoner
- |
  loneliness
- |
  lonely
- |
  loner
- |
  lonesome
- |
  lonesomely
- |
  lonesomeness
- |
  longboat
- |
  longbow
- |
  longevity
- |
  Longfellow
- |
  longhair
- |
  longhaired
- |
  longhand
- |
  longhorn
- |
  longhouse
- |
  longing
- |
  longingly
- |
  longish
- |
  longitude
- |
  longitudinal
- |
  longshore
- |
  longshoreman
- |
  longstanding
- |
  longtime
- |
  Longueuil
- |
  longueur
- |
  Lonna
- |
  Lonnie
- |
  Lonny
- |
  loofa
- |
  loofah
- |
  lookalike
- |
  looker
- |
  lookout
- |
  looks
- |
  looney
- |
  looniness
- |
  loony
- |
  looper
- |
  loophole
- |
  loopy
- |
  loose
- |
  loosely
- |
  loosen
- |
  looseness
- |
  loosening
- |
  looter
- |
  looting
- |
  loper
- |
  lopsided
- |
  lopsidedly
- |
  lopsidedness
- |
  loquacious
- |
  loquaciously
- |
  loquacity
- |
  Loraine
- |
  lordliness
- |
  lordly
- |
  Lordship
- |
  lordship
- |
  Lorelei
- |
  Loren
- |
  Lorene
- |
  Lorenzo
- |
  Loretta
- |
  lorgnette
- |
  lorgnettes
- |
  Lorinda
- |
  loris
- |
  Lorna
- |
  Lorraine
- |
  lorry
- |
  loser
- |
  losses
- |
  Lothario
- |
  Lothian
- |
  lotion
- |
  Lotta
- |
  lottery
- |
  Lottie
- |
  lotto
- |
  Lotty
- |
  lotus
- |
  louche
- |
  loudhailer
- |
  loudish
- |
  loudly
- |
  loudmouth
- |
  loudmouthed
- |
  loudness
- |
  loudspeaker
- |
  Louie
- |
  Louis
- |
  Louisa
- |
  Louise
- |
  Louisiana
- |
  Louisianan
- |
  Louisianian
- |
  Louisville
- |
  Louisvillian
- |
  lounge
- |
  lounger
- |
  Lourdes
- |
  loury
- |
  louse
- |
  lousily
- |
  lousiness
- |
  lousy
- |
  loutish
- |
  loutishly
- |
  louver
- |
  louvered
- |
  Louvre
- |
  louvre
- |
  louvred
- |
  lovability
- |
  lovable
- |
  loveable
- |
  lovebird
- |
  lovechild
- |
  Lovelace
- |
  loveless
- |
  lovelily
- |
  loveliness
- |
  lovelorn
- |
  lovely
- |
  lovemaking
- |
  lover
- |
  loverly
- |
  lovers
- |
  lovesick
- |
  lovesickness
- |
  loving
- |
  lovingly
- |
  lowball
- |
  lowborn
- |
  lowboy
- |
  lowbred
- |
  lowbrow
- |
  lowdown
- |
  Lowell
- |
  Lower
- |
  lower
- |
  lowercase
- |
  lowering
- |
  loweringly
- |
  lowermost
- |
  lowery
- |
  lowish
- |
  lowland
- |
  lowlander
- |
  Lowlands
- |
  lowlife
- |
  lowliness
- |
  lowlives
- |
  lowly
- |
  lowness
- |
  loyal
- |
  loyalism
- |
  Loyalist
- |
  loyalist
- |
  loyally
- |
  loyalty
- |
  Loyang
- |
  Loyola
- |
  lozenge
- |
  Luanda
- |
  Luanne
- |
  lubber
- |
  lubberly
- |
  Lubbock
- |
  Lubeck
- |
  Lublin
- |
  lubricant
- |
  lubricate
- |
  lubrication
- |
  lubricator
- |
  lubricious
- |
  lubriciously
- |
  lubricity
- |
  lubricous
- |
  Lubumbashi
- |
  lucency
- |
  lucent
- |
  lucently
- |
  Lucerne
- |
  lucerne
- |
  Lucia
- |
  Lucian
- |
  lucid
- |
  lucidity
- |
  lucidly
- |
  lucidness
- |
  Lucifer
- |
  lucifer
- |
  Lucile
- |
  Lucille
- |
  Lucinda
- |
  Lucite
- |
  Lucius
- |
  luckily
- |
  luckiness
- |
  luckless
- |
  Lucknow
- |
  lucky
- |
  lucrative
- |
  lucratively
- |
  lucre
- |
  Lucretia
- |
  Lucretian
- |
  Lucretius
- |
  lucubrate
- |
  lucubration
- |
  lucubrations
- |
  lucubrator
- |
  Luddite
- |
  Ludhiana
- |
  ludic
- |
  ludicrous
- |
  ludicrously
- |
  Ludwig
- |
  Luella
- |
  Luftwaffe
- |
  Lugansk
- |
  luggage
- |
  lugger
- |
  lugsail
- |
  lugubrious
- |
  lugubriously
- |
  lukewarm
- |
  lukewarmly
- |
  lukewarmness
- |
  lullaby
- |
  lumbago
- |
  lumbar
- |
  lumber
- |
  lumberer
- |
  lumbering
- |
  lumberjack
- |
  lumberman
- |
  lumberyard
- |
  lumen
- |
  lumenal
- |
  lumina
- |
  luminal
- |
  luminance
- |
  luminaria
- |
  luminary
- |
  luminescence
- |
  luminescent
- |
  luminosity
- |
  luminous
- |
  luminously
- |
  luminousness
- |
  lummox
- |
  lumpectomy
- |
  lumpen
- |
  lumpily
- |
  lumpiness
- |
  lumpish
- |
  lumpishly
- |
  lumpishness
- |
  lumps
- |
  lumpy
- |
  lunacy
- |
  lunar
- |
  lunate
- |
  lunatic
- |
  lunch
- |
  luncheon
- |
  luncheonette
- |
  lunchroom
- |
  lunchtime
- |
  lunette
- |
  lunge
- |
  lunged
- |
  lunger
- |
  lungfish
- |
  lunkhead
- |
  lunula
- |
  lunulae
- |
  Luoyang
- |
  lupin
- |
  lupine
- |
  Lupus
- |
  lupus
- |
  lurch
- |
  lurchingly
- |
  lurdan
- |
  lurdane
- |
  lurid
- |
  luridly
- |
  luridness
- |
  Lusaka
- |
  luscious
- |
  lusciously
- |
  lusciousness
- |
  lushly
- |
  lushness
- |
  Lushun
- |
  luster
- |
  lusterless
- |
  lustful
- |
  lustfully
- |
  lustfulness
- |
  lustily
- |
  lustiness
- |
  lustra
- |
  lustral
- |
  lustrate
- |
  lustration
- |
  lustre
- |
  lustrous
- |
  lustrously
- |
  lustrousness
- |
  lustrum
- |
  lusty
- |
  lutanist
- |
  lutecium
- |
  lutenist
- |
  lutetium
- |
  Luther
- |
  Lutheran
- |
  Lutheranism
- |
  lutist
- |
  Luton
- |
  luxate
- |
  luxation
- |
  Luxembourg
- |
  Luxembourger
- |
  Luxemburg
- |
  luxuriance
- |
  luxuriant
- |
  luxuriantly
- |
  luxuriate
- |
  luxuriation
- |
  luxurious
- |
  luxuriously
- |
  luxury
- |
  Luzon
- |
  Lyallpur
- |
  lycanthropic
- |
  lycanthropy
- |
  Lyceum
- |
  lyceum
- |
  lychee
- |
  Lycia
- |
  Lycian
- |
  Lycra
- |
  Lycurgus
- |
  Lydia
- |
  Lydian
- |
  Lyell
- |
  lying
- |
  Lyman
- |
  lymph
- |
  lymphatic
- |
  lymphocyte
- |
  lymphoid
- |
  lymphoma
- |
  lymphomata
- |
  lymphous
- |
  lynch
- |
  lyncher
- |
  lynching
- |
  lynchpin
- |
  Lynda
- |
  Lynette
- |
  Lynne
- |
  lyonnaise
- |
  Lyons
- |
  lyric
- |
  lyrical
- |
  lyrically
- |
  lyricism
- |
  lyricist
- |
  lyrics
- |
  lyses
- |
  lysin
- |
  lysis
- |
  Lysistrata
- |
  Maastricht
- |
  Mabel
- |
  macabre
- |
  macadam
- |
  macadamia
- |
  macadamize
- |
  Macanese
- |
  Macao
- |
  macaque
- |
  macarena
- |
  macaroni
- |
  macaronic
- |
  macaronics
- |
  macaroon
- |
  MacArthur
- |
  Macau
- |
  Macaulay
- |
  macaw
- |
  Macbeth
- |
  Maccabean
- |
  Maccabees
- |
  Maccabeus
- |
  MacDonald
- |
  Macdonald
- |
  Macedonia
- |
  Macedonian
- |
  macerate
- |
  maceration
- |
  macerator
- |
  machete
- |
  Machiavelli
- |
  machinable
- |
  machinate
- |
  machination
- |
  machinations
- |
  machinator
- |
  machine
- |
  machinery
- |
  machining
- |
  machinist
- |
  machismo
- |
  macho
- |
  macintosh
- |
  Mackenzie
- |
  mackerel
- |
  Mackinaw
- |
  mackinaw
- |
  mackintosh
- |
  MacLeish
- |
  Macmillan
- |
  Macon
- |
  macrame
- |
  macro
- |
  macrobiotic
- |
  macrobiotics
- |
  macrocephaly
- |
  macrocosm
- |
  macrocosmic
- |
  macrocosmos
- |
  macron
- |
  macrophage
- |
  macroscopic
- |
  Madagascan
- |
  Madagascar
- |
  Madam
- |
  madam
- |
  Madame
- |
  madame
- |
  madcap
- |
  madden
- |
  maddening
- |
  maddeningly
- |
  madder
- |
  madding
- |
  Madeira
- |
  Madeiran
- |
  Madeleine
- |
  Madeline
- |
  Madelyn
- |
  Mademoiselle
- |
  mademoiselle
- |
  Madge
- |
  madhouse
- |
  Madison
- |
  Madisonian
- |
  madly
- |
  madman
- |
  madness
- |
  Madonna
- |
  Madras
- |
  madras
- |
  Madrid
- |
  madrigal
- |
  madrigalian
- |
  madrigalist
- |
  Madrilenian
- |
  madrona
- |
  madrone
- |
  madrono
- |
  Madura
- |
  Madurai
- |
  madwoman
- |
  maelstrom
- |
  maenad
- |
  maenadic
- |
  maestoso
- |
  maestri
- |
  maestro
- |
  Maeterlinck
- |
  Mafia
- |
  mafia
- |
  Mafiosi
- |
  mafiosi
- |
  Mafioso
- |
  mafioso
- |
  magazine
- |
  Magdalena
- |
  Magdalene
- |
  Magdeburg
- |
  Magellan
- |
  magenta
- |
  Maggie
- |
  maggot
- |
  maggoty
- |
  Magherafelt
- |
  magic
- |
  magical
- |
  magically
- |
  magician
- |
  magisterial
- |
  magistracy
- |
  magistral
- |
  magistrate
- |
  magma
- |
  magmata
- |
  magmatic
- |
  magnanimity
- |
  magnanimous
- |
  magnate
- |
  magnesia
- |
  magnesium
- |
  magnet
- |
  magnetic
- |
  magnetically
- |
  magnetise
- |
  magnetism
- |
  magnetite
- |
  magnetizable
- |
  magnetize
- |
  magnetizer
- |
  magneto
- |
  magnetometer
- |
  magnifiable
- |
  magnificence
- |
  magnificent
- |
  magnifier
- |
  magnify
- |
  magniloquent
- |
  Magnitogorsk
- |
  magnitude
- |
  magnolia
- |
  magnum
- |
  magpie
- |
  Magritte
- |
  maguey
- |
  Magus
- |
  magus
- |
  Magyar
- |
  maharaja
- |
  maharajah
- |
  maharanee
- |
  maharani
- |
  maharishi
- |
  Mahatma
- |
  mahatma
- |
  Mahayana
- |
  Mahdi
- |
  Mahdism
- |
  Mahdist
- |
  Mahfouz
- |
  Mahican
- |
  mahjong
- |
  mahjongg
- |
  Mahler
- |
  mahogany
- |
  Mahomet
- |
  mahout
- |
  maiden
- |
  maidenhair
- |
  maidenhead
- |
  maidenhood
- |
  maidenly
- |
  maidservant
- |
  Maidstone
- |
  Maidu
- |
  maieutic
- |
  mailbag
- |
  mailbox
- |
  mailed
- |
  Mailer
- |
  mailer
- |
  mailing
- |
  Maillol
- |
  maillot
- |
  mailman
- |
  mails
- |
  mailwoman
- |
  maimer
- |
  Maimonides
- |
  Maine
- |
  Mainer
- |
  mainframe
- |
  mainland
- |
  mainline
- |
  mainliner
- |
  mainly
- |
  mainmast
- |
  mainsail
- |
  mainspring
- |
  mainstay
- |
  mainstream
- |
  maintain
- |
  maintainable
- |
  maintenance
- |
  maintop
- |
  Mainz
- |
  maiolica
- |
  maisonette
- |
  maize
- |
  majestic
- |
  majestically
- |
  Majesty
- |
  majesty
- |
  majolica
- |
  Major
- |
  major
- |
  Majorca
- |
  Majorcan
- |
  majordomo
- |
  majorette
- |
  majority
- |
  majorly
- |
  Majuro
- |
  majuscular
- |
  majuscule
- |
  Makalu
- |
  Makarios
- |
  makeover
- |
  maker
- |
  makeshift
- |
  makeup
- |
  making
- |
  makings
- |
  Makiyivka
- |
  makuta
- |
  Malabar
- |
  Malabo
- |
  Malacca
- |
  Malachi
- |
  Malachias
- |
  malachite
- |
  maladapted
- |
  maladjusted
- |
  maladroit
- |
  maladroitly
- |
  malady
- |
  Malaga
- |
  Malagasy
- |
  malaise
- |
  Malamud
- |
  malamute
- |
  Malang
- |
  malapert
- |
  Malaprop
- |
  malaprop
- |
  malapropism
- |
  malapropos
- |
  malaria
- |
  malarial
- |
  malarkey
- |
  malarky
- |
  Malathion
- |
  malathion
- |
  Malatya
- |
  Malawi
- |
  Malawian
- |
  Malay
- |
  Malaya
- |
  Malayalam
- |
  Malayan
- |
  Malaysia
- |
  Malaysian
- |
  Malcolm
- |
  malcontent
- |
  malcontented
- |
  Maldivan
- |
  Maldives
- |
  Maldivian
- |
  Malecite
- |
  malediction
- |
  maledictive
- |
  maledictory
- |
  malefaction
- |
  malefactor
- |
  malefic
- |
  maleficence
- |
  maleficent
- |
  maleness
- |
  malevolence
- |
  malevolent
- |
  malevolently
- |
  malfeasance
- |
  malfeasant
- |
  malformation
- |
  malformed
- |
  malfunction
- |
  Malian
- |
  malice
- |
  malicious
- |
  maliciously
- |
  malign
- |
  malignancy
- |
  malignant
- |
  malignantly
- |
  maligner
- |
  malignity
- |
  malignly
- |
  malinger
- |
  malingerer
- |
  Malinowski
- |
  Maliseet
- |
  malison
- |
  mallard
- |
  Mallarme
- |
  malleability
- |
  malleable
- |
  malleably
- |
  mallei
- |
  mallet
- |
  malleus
- |
  Mallory
- |
  mallow
- |
  Malmo
- |
  malmsey
- |
  malnourished
- |
  malnutrition
- |
  malocclusion
- |
  malodor
- |
  malodorous
- |
  malodorously
- |
  Malory
- |
  maloti
- |
  malpractice
- |
  Malraux
- |
  Malta
- |
  malted
- |
  Maltese
- |
  Malthus
- |
  Malthusian
- |
  maltose
- |
  maltreat
- |
  maltreatment
- |
  malty
- |
  malversation
- |
  Malvinas
- |
  mamba
- |
  mambo
- |
  Mamet
- |
  Mamie
- |
  mamma
- |
  mammal
- |
  mammalian
- |
  mammalogist
- |
  mammalogy
- |
  mammary
- |
  mammogram
- |
  mammography
- |
  Mammon
- |
  mammon
- |
  mammonism
- |
  mammonist
- |
  mammoth
- |
  mammy
- |
  Mamore
- |
  manacle
- |
  manacles
- |
  manage
- |
  manageable
- |
  manageably
- |
  management
- |
  manager
- |
  managerial
- |
  managerially
- |
  managership
- |
  Managua
- |
  Managuan
- |
  Manama
- |
  manana
- |
  Manaos
- |
  manat
- |
  manatee
- |
  Manaus
- |
  Manchester
- |
  Manchu
- |
  Manchuria
- |
  Manchurian
- |
  manciple
- |
  Mancunian
- |
  mandala
- |
  Mandalay
- |
  mandalic
- |
  mandamus
- |
  Mandan
- |
  Mandarin
- |
  mandarin
- |
  mandarinate
- |
  mandarinism
- |
  mandate
- |
  mandatorily
- |
  mandatory
- |
  Mandela
- |
  Mandelstam
- |
  mandible
- |
  mandibular
- |
  mandibulate
- |
  Mandingo
- |
  mandolin
- |
  mandolinist
- |
  mandrake
- |
  mandrel
- |
  mandril
- |
  mandrill
- |
  Mandy
- |
  maned
- |
  manege
- |
  Manes
- |
  manes
- |
  Manet
- |
  maneuver
- |
  maneuverable
- |
  maneuvering
- |
  maneuvers
- |
  Manfred
- |
  manful
- |
  manfully
- |
  manfulness
- |
  manganese
- |
  mange
- |
  manger
- |
  mangily
- |
  manginess
- |
  mangle
- |
  mangler
- |
  mango
- |
  mangrove
- |
  mangy
- |
  manhandle
- |
  Manhattan
- |
  manhattan
- |
  Manhattanite
- |
  manhole
- |
  manhood
- |
  manhunt
- |
  mania
- |
  maniac
- |
  maniacal
- |
  maniacally
- |
  manic
- |
  manically
- |
  Manichaeism
- |
  Manicheism
- |
  manicotti
- |
  manicure
- |
  manicurist
- |
  manifest
- |
  manifestly
- |
  manifesto
- |
  manifold
- |
  manifoldly
- |
  manifoldness
- |
  manikin
- |
  Manila
- |
  manioc
- |
  manipulable
- |
  manipulate
- |
  manipulation
- |
  manipulative
- |
  manipulator
- |
  manipulatory
- |
  Manitoba
- |
  Manitoban
- |
  manitou
- |
  Manitoulin
- |
  Manizales
- |
  mankind
- |
  Manley
- |
  manlike
- |
  manliness
- |
  manly
- |
  manmade
- |
  manna
- |
  manned
- |
  mannequin
- |
  manner
- |
  mannered
- |
  mannerism
- |
  mannerist
- |
  mannerliness
- |
  mannerly
- |
  manners
- |
  Mannheim
- |
  mannikin
- |
  mannish
- |
  mannishly
- |
  mannishness
- |
  manoeuvre
- |
  manoeuvring
- |
  manometer
- |
  manometric
- |
  manometrical
- |
  manometry
- |
  manor
- |
  manorial
- |
  manorialism
- |
  manpower
- |
  manque
- |
  mansard
- |
  manse
- |
  manservant
- |
  mansion
- |
  manslaughter
- |
  manslayer
- |
  mansuetude
- |
  manta
- |
  manteau
- |
  Mantegna
- |
  mantel
- |
  mantelpiece
- |
  mantes
- |
  mantic
- |
  mantilla
- |
  mantis
- |
  mantissa
- |
  mantle
- |
  mantra
- |
  mantric
- |
  Mantua
- |
  manual
- |
  manually
- |
  Manuel
- |
  manufactory
- |
  manufacture
- |
  manufacturer
- |
  manumission
- |
  manumit
- |
  manumitter
- |
  manure
- |
  manurial
- |
  manuscript
- |
  Manxman
- |
  Manxwoman
- |
  manyfold
- |
  manzanita
- |
  Maoism
- |
  Maoist
- |
  Maori
- |
  maple
- |
  mapmaker
- |
  mappable
- |
  mapper
- |
  Maputo
- |
  maquiladora
- |
  maquis
- |
  marabou
- |
  maraca
- |
  Maracaibo
- |
  Maracay
- |
  Maranon
- |
  maraschino
- |
  Marat
- |
  Marathi
- |
  Marathon
- |
  marathon
- |
  marathoner
- |
  marathoning
- |
  maraud
- |
  marauder
- |
  marauding
- |
  marble
- |
  marbled
- |
  marbleize
- |
  marbles
- |
  marbling
- |
  marbly
- |
  marcasite
- |
  Marcel
- |
  marcel
- |
  Marcella
- |
  Marcellus
- |
  March
- |
  march
- |
  marcher
- |
  marchioness
- |
  Marcia
- |
  Marciano
- |
  Marconi
- |
  Marcos
- |
  Marcus
- |
  Marcuse
- |
  Margaret
- |
  margarine
- |
  margarita
- |
  Margery
- |
  Margie
- |
  margin
- |
  marginal
- |
  marginalia
- |
  marginalise
- |
  marginalize
- |
  marginally
- |
  Margo
- |
  Margot
- |
  margrave
- |
  Margrethe
- |
  Marguerite
- |
  marguerite
- |
  Maria
- |
  maria
- |
  mariachi
- |
  Marian
- |
  Mariana
- |
  Marianas
- |
  Marianna
- |
  Marianne
- |
  maricultural
- |
  mariculture
- |
  Marie
- |
  Marietta
- |
  marigold
- |
  marihuana
- |
  marijuana
- |
  Marilee
- |
  Marilyn
- |
  Marilynn
- |
  marimba
- |
  Marin
- |
  Marina
- |
  marina
- |
  marinade
- |
  marinara
- |
  marinate
- |
  marination
- |
  Marinduque
- |
  Marine
- |
  marine
- |
  mariner
- |
  Marines
- |
  Mario
- |
  Mariolatry
- |
  Marion
- |
  marionette
- |
  marital
- |
  maritally
- |
  maritime
- |
  Maritimer
- |
  Mariupol
- |
  Marius
- |
  marjoram
- |
  Marjorie
- |
  Marjory
- |
  marka
- |
  Markab
- |
  markdown
- |
  marked
- |
  markedly
- |
  marker
- |
  market
- |
  marketable
- |
  marketeer
- |
  marketer
- |
  marketing
- |
  marketplace
- |
  Markham
- |
  marking
- |
  markka
- |
  markkaa
- |
  marks
- |
  marksman
- |
  marksmanship
- |
  markswoman
- |
  markup
- |
  Marla
- |
  Marlborough
- |
  Marlene
- |
  Marlin
- |
  marlin
- |
  marlinespike
- |
  marlinspike
- |
  Marlowe
- |
  marly
- |
  Marlyn
- |
  marmalade
- |
  Marmara
- |
  marmoreal
- |
  marmoset
- |
  marmot
- |
  Marne
- |
  maroon
- |
  Marquand
- |
  marque
- |
  marquee
- |
  Marquesan
- |
  Marquesas
- |
  marquess
- |
  marqueterie
- |
  marquetery
- |
  marquetry
- |
  Marquette
- |
  marquis
- |
  marquise
- |
  marquisette
- |
  Marrakech
- |
  Marrakesh
- |
  marriage
- |
  marriageable
- |
  married
- |
  marrow
- |
  marrowbone
- |
  marry
- |
  Marseille
- |
  Marseilles
- |
  marsh
- |
  Marsha
- |
  Marshal
- |
  marshal
- |
  marshaler
- |
  Marshall
- |
  marshalship
- |
  marshiness
- |
  marshmallow
- |
  marshy
- |
  marsupial
- |
  Marta
- |
  Martel
- |
  marten
- |
  Martha
- |
  Marti
- |
  Martial
- |
  martial
- |
  martially
- |
  Martian
- |
  martian
- |
  Martin
- |
  martin
- |
  martinet
- |
  martingale
- |
  martini
- |
  Martinique
- |
  martyr
- |
  martyrdom
- |
  martyrize
- |
  Marva
- |
  marvel
- |
  Marvell
- |
  marvellous
- |
  marvellously
- |
  marvelous
- |
  marvelously
- |
  Marvin
- |
  Marxian
- |
  Marxism
- |
  Marxist
- |
  Maryann
- |
  Maryanne
- |
  Maryellen
- |
  Maryland
- |
  Marylander
- |
  Marylon
- |
  Marylyn
- |
  marzipan
- |
  Masai
- |
  Masaryk
- |
  Masbate
- |
  mascara
- |
  mascot
- |
  masculine
- |
  masculinely
- |
  masculinity
- |
  Masefield
- |
  maser
- |
  Maseru
- |
  masher
- |
  Mashhad
- |
  masked
- |
  masker
- |
  masochism
- |
  masochist
- |
  masochistic
- |
  Mason
- |
  mason
- |
  Masonic
- |
  Masonry
- |
  masonry
- |
  masque
- |
  masquer
- |
  masquerade
- |
  masquerader
- |
  Massachuset
- |
  Massachusett
- |
  massacre
- |
  massage
- |
  Massasoit
- |
  Massenet
- |
  masses
- |
  masseur
- |
  masseuse
- |
  massif
- |
  Massilia
- |
  massive
- |
  massively
- |
  massiveness
- |
  massless
- |
  massy
- |
  mastectomy
- |
  masted
- |
  Master
- |
  master
- |
  masterful
- |
  masterfully
- |
  masterliness
- |
  masterly
- |
  mastermind
- |
  masterpiece
- |
  Masters
- |
  masterstroke
- |
  masterwork
- |
  mastery
- |
  masthead
- |
  mastic
- |
  masticate
- |
  mastication
- |
  masticator
- |
  masticatory
- |
  mastiff
- |
  mastitis
- |
  mastodon
- |
  mastoid
- |
  masturbate
- |
  masturbation
- |
  masturbator
- |
  masturbatory
- |
  Matabeleland
- |
  matador
- |
  Matamoros
- |
  match
- |
  matchbook
- |
  matchbox
- |
  matched
- |
  matcher
- |
  matching
- |
  matchless
- |
  matchlock
- |
  matchmaker
- |
  matchmaking
- |
  matchstick
- |
  matchup
- |
  matchwood
- |
  material
- |
  materialise
- |
  materialism
- |
  materialist
- |
  materialize
- |
  materially
- |
  materials
- |
  materiel
- |
  maternal
- |
  maternalism
- |
  maternalist
- |
  maternally
- |
  maternity
- |
  mathematic
- |
  mathematical
- |
  mathematics
- |
  Mather
- |
  Mathilda
- |
  maths
- |
  matinee
- |
  matins
- |
  Matisse
- |
  Matlock
- |
  matriarch
- |
  matriarchal
- |
  matriarchic
- |
  matriarchy
- |
  matrices
- |
  matricidal
- |
  matricide
- |
  matriculant
- |
  matriculate
- |
  matrilineal
- |
  matrimonial
- |
  matrimony
- |
  matrix
- |
  matron
- |
  matronhood
- |
  matronliness
- |
  matronly
- |
  Matsu
- |
  matte
- |
  matted
- |
  matter
- |
  Matterhorn
- |
  Matthew
- |
  Matthias
- |
  matting
- |
  mattins
- |
  mattock
- |
  mattress
- |
  maturate
- |
  maturation
- |
  maturational
- |
  mature
- |
  maturely
- |
  matureness
- |
  maturity
- |
  matutinal
- |
  matzo
- |
  matzoh
- |
  matzot
- |
  matzoth
- |
  Maude
- |
  maudlin
- |
  Maugham
- |
  mauler
- |
  maunder
- |
  Maupassant
- |
  Maureen
- |
  Mauretania
- |
  Mauretanian
- |
  Mauriac
- |
  Maurice
- |
  Maurine
- |
  Mauritania
- |
  Mauritanian
- |
  Mauritian
- |
  Mauritius
- |
  Maurois
- |
  mausolea
- |
  mausoleum
- |
  mauve
- |
  mauvish
- |
  maven
- |
  maverick
- |
  mavin
- |
  mawkish
- |
  mawkishly
- |
  mawkishness
- |
  maxilla
- |
  maxillae
- |
  maxillary
- |
  maxim
- |
  maxima
- |
  maximal
- |
  maximally
- |
  Maximilian
- |
  maximise
- |
  maximization
- |
  maximize
- |
  maximizer
- |
  maximum
- |
  Maxine
- |
  Maxwell
- |
  Mayaguez
- |
  Mayan
- |
  mayapple
- |
  maybe
- |
  Mayday
- |
  mayday
- |
  mayflower
- |
  mayfly
- |
  mayhem
- |
  Maynard
- |
  mayonnaise
- |
  mayor
- |
  mayoral
- |
  mayoralty
- |
  mayoress
- |
  mayorship
- |
  Maypole
- |
  maypole
- |
  Mazarin
- |
  Mazatlan
- |
  mazourka
- |
  mazurka
- |
  Mazzini
- |
  Mbabane
- |
  Mbini
- |
  Mboya
- |
  McAllen
- |
  McCarthy
- |
  McCarthyism
- |
  McCartney
- |
  McClellan
- |
  McCormick
- |
  McCoy
- |
  McCullers
- |
  McGovern
- |
  McGuffey
- |
  McJob
- |
  McKinley
- |
  McLuhan
- |
  Meade
- |
  meadow
- |
  meadowland
- |
  meadowlark
- |
  meadowsweet
- |
  meadowy
- |
  meager
- |
  meagerly
- |
  meagerness
- |
  meagre
- |
  mealiness
- |
  mealtime
- |
  mealy
- |
  mealybug
- |
  mealymouthed
- |
  meander
- |
  meandering
- |
  meanderings
- |
  meanders
- |
  meandrous
- |
  meanie
- |
  meaning
- |
  meaningful
- |
  meaningfully
- |
  meaningless
- |
  meaningly
- |
  meanly
- |
  meanness
- |
  means
- |
  meant
- |
  meantime
- |
  meanwhile
- |
  Meany
- |
  meany
- |
  measles
- |
  measly
- |
  measurable
- |
  measurably
- |
  measure
- |
  measured
- |
  measureless
- |
  measurement
- |
  measurer
- |
  measures
- |
  meatball
- |
  meatiness
- |
  meatless
- |
  meatloaf
- |
  meatpacking
- |
  meaty
- |
  Mecca
- |
  mecca
- |
  mechanic
- |
  mechanical
- |
  mechanically
- |
  mechanics
- |
  mechanise
- |
  mechanism
- |
  mechanistic
- |
  mechanize
- |
  mechanized
- |
  mechanizer
- |
  medal
- |
  medalist
- |
  medallion
- |
  medallist
- |
  Medan
- |
  meddle
- |
  meddler
- |
  meddlesome
- |
  Medea
- |
  Medellin
- |
  medevac
- |
  Media
- |
  media
- |
  mediacy
- |
  mediaeval
- |
  medial
- |
  medially
- |
  Median
- |
  median
- |
  medianly
- |
  mediate
- |
  mediately
- |
  mediation
- |
  mediator
- |
  mediatory
- |
  medic
- |
  medicable
- |
  Medicaid
- |
  medicaid
- |
  medical
- |
  medically
- |
  medicament
- |
  Medicare
- |
  medicare
- |
  medicate
- |
  medicated
- |
  medication
- |
  medicative
- |
  Medicean
- |
  Medici
- |
  medicinal
- |
  medicinally
- |
  medicine
- |
  medico
- |
  medieval
- |
  medievalism
- |
  medievalist
- |
  medievally
- |
  Medigap
- |
  Medina
- |
  mediocre
- |
  mediocrely
- |
  mediocrity
- |
  meditate
- |
  meditation
- |
  meditational
- |
  meditative
- |
  meditatively
- |
  meditator
- |
  medium
- |
  mediumism
- |
  mediumistic
- |
  mediumship
- |
  medley
- |
  medulla
- |
  medullae
- |
  medullar
- |
  medullary
- |
  Medusa
- |
  medusa
- |
  meekly
- |
  meekness
- |
  meerkat
- |
  meerschaum
- |
  Meerut
- |
  meeting
- |
  meetinghouse
- |
  meetly
- |
  megabit
- |
  megabuck
- |
  megabyte
- |
  megacycle
- |
  megadeath
- |
  megadose
- |
  megafauna
- |
  megaflops
- |
  megahertz
- |
  megalith
- |
  Megalithic
- |
  megalithic
- |
  megalomania
- |
  megalomaniac
- |
  megalomanic
- |
  megalopolis
- |
  Megan
- |
  megaphone
- |
  megaton
- |
  megatonnage
- |
  megavitamin
- |
  megawatt
- |
  megawattage
- |
  Megillah
- |
  Megrez
- |
  megrim
- |
  meioses
- |
  meiosis
- |
  meiotic
- |
  meiotically
- |
  meitnerium
- |
  Meknes
- |
  Mekong
- |
  melamine
- |
  melancholia
- |
  melancholiac
- |
  melancholic
- |
  melancholy
- |
  Melanesia
- |
  Melanesian
- |
  melange
- |
  melanic
- |
  Melanie
- |
  melanin
- |
  melanism
- |
  melanistic
- |
  melanoma
- |
  melanomata
- |
  melanosis
- |
  melanotic
- |
  melatonin
- |
  Melba
- |
  Melbourne
- |
  melee
- |
  Melian
- |
  Melinda
- |
  meliorable
- |
  meliorate
- |
  melioration
- |
  meliorative
- |
  meliorism
- |
  meliorist
- |
  melioristic
- |
  Melissa
- |
  mellifluence
- |
  mellifluent
- |
  mellifluous
- |
  Mellon
- |
  mellow
- |
  mellowly
- |
  mellowness
- |
  melodeon
- |
  melodic
- |
  melodically
- |
  melodious
- |
  melodiously
- |
  melodrama
- |
  melodramatic
- |
  melody
- |
  melon
- |
  Melos
- |
  meltable
- |
  meltdown
- |
  meltingly
- |
  meltwater
- |
  Melva
- |
  Melville
- |
  Melvillean
- |
  Melvin
- |
  Melvyn
- |
  member
- |
  membership
- |
  membranal
- |
  membrane
- |
  membraneous
- |
  membranous
- |
  memento
- |
  memetic
- |
  Memling
- |
  memoir
- |
  memoirist
- |
  memoirs
- |
  memorabilia
- |
  memorability
- |
  memorable
- |
  memorably
- |
  memoranda
- |
  memorandum
- |
  memorial
- |
  memorialize
- |
  memorially
- |
  memorise
- |
  memorization
- |
  memorize
- |
  memorizer
- |
  memory
- |
  Memphis
- |
  memsahib
- |
  menace
- |
  menacer
- |
  menacing
- |
  menacingly
- |
  menage
- |
  menagerie
- |
  Menander
- |
  menarche
- |
  menarcheal
- |
  Mencius
- |
  Mencken
- |
  mendable
- |
  mendacious
- |
  mendaciously
- |
  mendacity
- |
  Mendel
- |
  Mendeleev
- |
  mendelevium
- |
  Mendelian
- |
  Mendelssohn
- |
  mender
- |
  mendicancy
- |
  mendicant
- |
  Menelaus
- |
  Menes
- |
  menfolk
- |
  menfolks
- |
  Mengzi
- |
  menhaden
- |
  menhir
- |
  menial
- |
  menially
- |
  meningeal
- |
  meninges
- |
  meningitis
- |
  meninx
- |
  menisci
- |
  meniscoid
- |
  meniscus
- |
  Menkar
- |
  Mennonite
- |
  menopausal
- |
  menopause
- |
  Menorah
- |
  menorah
- |
  Menotti
- |
  Mensa
- |
  mensch
- |
  menschen
- |
  menservants
- |
  menses
- |
  menstrual
- |
  menstruate
- |
  menstruation
- |
  mensurable
- |
  mensural
- |
  mensuration
- |
  menswear
- |
  mental
- |
  mentalist
- |
  mentality
- |
  mentally
- |
  mentation
- |
  menthol
- |
  mentholated
- |
  mention
- |
  mentionable
- |
  mentor
- |
  mentorship
- |
  mephitic
- |
  mephitical
- |
  mephitis
- |
  Merak
- |
  mercantile
- |
  mercantilism
- |
  mercantilist
- |
  Mercator
- |
  mercenarily
- |
  mercenary
- |
  mercer
- |
  mercerize
- |
  merchandise
- |
  merchandiser
- |
  merchandize
- |
  merchandizer
- |
  merchant
- |
  merchantable
- |
  merchantman
- |
  Mercia
- |
  Mercian
- |
  merciful
- |
  mercifully
- |
  mercifulness
- |
  merciless
- |
  mercilessly
- |
  mercurial
- |
  mercuriality
- |
  mercurially
- |
  mercuric
- |
  mercurous
- |
  Mercury
- |
  mercury
- |
  mercy
- |
  Meredith
- |
  merely
- |
  merengue
- |
  meretricious
- |
  merganser
- |
  merge
- |
  merger
- |
  Merida
- |
  meridian
- |
  meringue
- |
  merino
- |
  merit
- |
  meritless
- |
  meritocracy
- |
  meritocrat
- |
  meritocratic
- |
  meritorious
- |
  merits
- |
  Merle
- |
  Merlin
- |
  Merlyn
- |
  mermaid
- |
  merman
- |
  meronym
- |
  meronymous
- |
  meronymy
- |
  Merrill
- |
  Merrily
- |
  merrily
- |
  merriment
- |
  merriness
- |
  Merry
- |
  merry
- |
  merrymaker
- |
  merrymaking
- |
  Mersey
- |
  Merseyside
- |
  Mersin
- |
  Merton
- |
  Mervin
- |
  Mervyn
- |
  Merwin
- |
  Merwyn
- |
  mesalliance
- |
  mescal
- |
  mescaline
- |
  mesclun
- |
  Mesdames
- |
  mesdames
- |
  Meshed
- |
  meshed
- |
  meshes
- |
  meshuga
- |
  meshugaas
- |
  meshugah
- |
  meshugga
- |
  meshuggener
- |
  meshwork
- |
  mesial
- |
  mesmeric
- |
  mesmerise
- |
  mesmerism
- |
  mesmerist
- |
  mesmerize
- |
  mesmerized
- |
  mesmerizer
- |
  mesmerizing
- |
  mesne
- |
  Mesoamerica
- |
  Mesoamerican
- |
  Mesolithic
- |
  mesomorph
- |
  mesomorphic
- |
  meson
- |
  Mesopotamia
- |
  Mesopotamian
- |
  mesosphere
- |
  mesospheric
- |
  Mesozoic
- |
  mesquit
- |
  Mesquite
- |
  mesquite
- |
  message
- |
  messeigneurs
- |
  messenger
- |
  Messiah
- |
  messiah
- |
  messiahship
- |
  Messianic
- |
  messianic
- |
  Messianism
- |
  Messias
- |
  Messieurs
- |
  messieurs
- |
  messily
- |
  Messina
- |
  messiness
- |
  messmate
- |
  messy
- |
  mestiza
- |
  mestizo
- |
  metabolic
- |
  metabolism
- |
  metabolite
- |
  metabolize
- |
  metacarpal
- |
  metacarpi
- |
  metacarpus
- |
  Metacom
- |
  metafiction
- |
  Metairie
- |
  metal
- |
  metalanguage
- |
  metallic
- |
  metallically
- |
  metallurgic
- |
  metallurgist
- |
  metallurgy
- |
  metalware
- |
  metalwork
- |
  metalworker
- |
  metalworking
- |
  metamorphic
- |
  metamorphism
- |
  metamorphose
- |
  metamorphous
- |
  metanoia
- |
  metaphor
- |
  metaphoric
- |
  metaphorical
- |
  metaphysical
- |
  metaphysics
- |
  metastases
- |
  metastasis
- |
  metastasize
- |
  metastatic
- |
  metatarsal
- |
  metatarsi
- |
  metatarsus
- |
  metatheses
- |
  metathesis
- |
  metathesize
- |
  metathetic
- |
  metathetical
- |
  meteor
- |
  meteoric
- |
  meteorically
- |
  meteorite
- |
  meteoritic
- |
  meteoritical
- |
  meteoroid
- |
  meteorologic
- |
  meteorology
- |
  meter
- |
  meterage
- |
  methadon
- |
  methadone
- |
  methane
- |
  methanol
- |
  methaqualone
- |
  methinks
- |
  method
- |
  methodic
- |
  methodical
- |
  methodically
- |
  Methodism
- |
  Methodist
- |
  Methodistic
- |
  methodize
- |
  methodology
- |
  methought
- |
  Methuselah
- |
  methyl
- |
  methylic
- |
  metical
- |
  meticulosity
- |
  meticulous
- |
  meticulously
- |
  metier
- |
  Metis
- |
  metis
- |
  metonym
- |
  metonymic
- |
  metonymical
- |
  metonymy
- |
  metre
- |
  metric
- |
  metrical
- |
  metrically
- |
  metricate
- |
  metrication
- |
  metricize
- |
  metrics
- |
  Metro
- |
  metro
- |
  metronome
- |
  metronomic
- |
  metroplex
- |
  metropolis
- |
  metropolitan
- |
  Metternich
- |
  mettle
- |
  mettlesome
- |
  Meuse
- |
  Mexicali
- |
  Mexican
- |
  Mexico
- |
  Meyerbeer
- |
  mezuza
- |
  mezuzah
- |
  mezuzot
- |
  mezuzoth
- |
  mezzanine
- |
  mezzo
- |
  mezzotint
- |
  mezzotinter
- |
  Miami
- |
  Miamian
- |
  miasma
- |
  miasmal
- |
  miasmata
- |
  miasmatic
- |
  miasmic
- |
  miasmically
- |
  Micah
- |
  Michael
- |
  Micheas
- |
  Michelangelo
- |
  Michele
- |
  Michelle
- |
  Michigan
- |
  Michigander
- |
  Michiganite
- |
  Michoacan
- |
  Mickey
- |
  mickey
- |
  Micmac
- |
  micra
- |
  micro
- |
  microbe
- |
  microbial
- |
  microbic
- |
  microbiology
- |
  microbrew
- |
  microbrewer
- |
  microbrewery
- |
  microburst
- |
  microbus
- |
  microcapsule
- |
  microcephaly
- |
  microchip
- |
  microcircuit
- |
  microcosm
- |
  microcosmic
- |
  microcosmos
- |
  microdot
- |
  microfiber
- |
  microfiche
- |
  microfilm
- |
  microfloppy
- |
  micrograph
- |
  microgroove
- |
  microlight
- |
  microlith
- |
  microlithic
- |
  micromanage
- |
  micromanager
- |
  micrometer
- |
  micron
- |
  Micronesia
- |
  Micronesian
- |
  microphone
- |
  microscope
- |
  microscopic
- |
  Microscopium
- |
  microscopy
- |
  microsecond
- |
  microsurgery
- |
  microwavable
- |
  microwave
- |
  micturate
- |
  micturition
- |
  midair
- |
  Midas
- |
  midday
- |
  midden
- |
  middle
- |
  middlebrow
- |
  middleman
- |
  middlemost
- |
  middleweight
- |
  middling
- |
  middlingly
- |
  middy
- |
  Mideast
- |
  Mideastern
- |
  Mideasterner
- |
  midge
- |
  midget
- |
  Midian
- |
  Midianite
- |
  Midland
- |
  midland
- |
  Midlands
- |
  midlife
- |
  midline
- |
  midmost
- |
  midnight
- |
  midpoint
- |
  midrib
- |
  midriff
- |
  midsection
- |
  midshipman
- |
  midships
- |
  midsize
- |
  midst
- |
  midstream
- |
  midsummer
- |
  midterm
- |
  midtown
- |
  Midway
- |
  midway
- |
  midweek
- |
  midweekly
- |
  Midwest
- |
  Midwestern
- |
  Midwesterner
- |
  midwife
- |
  midwifery
- |
  midwinter
- |
  midwives
- |
  midyear
- |
  miffed
- |
  miffy
- |
  might
- |
  mightily
- |
  mightiness
- |
  mighty
- |
  mignonette
- |
  migraine
- |
  migrainous
- |
  migrant
- |
  migrate
- |
  migration
- |
  migrational
- |
  migrator
- |
  migratory
- |
  mikado
- |
  mikva
- |
  mikvah
- |
  mikveh
- |
  mikvos
- |
  mikvot
- |
  mikvoth
- |
  miladi
- |
  milady
- |
  Milan
- |
  Milanese
- |
  milch
- |
  mildew
- |
  mildewy
- |
  mildish
- |
  mildly
- |
  mildness
- |
  Mildred
- |
  mileage
- |
  milepost
- |
  miler
- |
  Miles
- |
  milestone
- |
  Miletus
- |
  Milford
- |
  Milicent
- |
  milieu
- |
  milieux
- |
  militance
- |
  militancy
- |
  militant
- |
  militantly
- |
  militarily
- |
  militarism
- |
  militarist
- |
  militaristic
- |
  militarize
- |
  military
- |
  militate
- |
  militia
- |
  militiaman
- |
  milker
- |
  milkiness
- |
  milking
- |
  milkmaid
- |
  milkman
- |
  milkshake
- |
  milksop
- |
  milkweed
- |
  milky
- |
  millage
- |
  Millard
- |
  Millay
- |
  milldam
- |
  millenarian
- |
  millenary
- |
  millennia
- |
  millennial
- |
  millennially
- |
  millennium
- |
  millepede
- |
  Miller
- |
  miller
- |
  Millet
- |
  millet
- |
  milliampere
- |
  milliard
- |
  millibar
- |
  Millicent
- |
  Millie
- |
  milligram
- |
  milligramme
- |
  milliliter
- |
  millime
- |
  millimeter
- |
  millimetre
- |
  milliner
- |
  millinery
- |
  milling
- |
  million
- |
  millionaire
- |
  millionnaire
- |
  millionth
- |
  millipede
- |
  millisecond
- |
  millivolt
- |
  millpond
- |
  millrace
- |
  millstone
- |
  millstream
- |
  millwright
- |
  Milne
- |
  milord
- |
  Milosevic
- |
  Milosz
- |
  Milquetoast
- |
  milquetoast
- |
  Milton
- |
  Milwaukee
- |
  mimeograph
- |
  mimer
- |
  mimesis
- |
  mimetic
- |
  mimetically
- |
  mimic
- |
  mimicker
- |
  mimicry
- |
  mimosa
- |
  minable
- |
  minacious
- |
  minaret
- |
  minareted
- |
  minatorial
- |
  minatory
- |
  mince
- |
  mincemeat
- |
  mincer
- |
  mincing
- |
  mincingly
- |
  Mindanao
- |
  mindblower
- |
  minded
- |
  minder
- |
  mindful
- |
  mindfully
- |
  mindfulness
- |
  mindless
- |
  mindlessly
- |
  mindlessness
- |
  Mindoro
- |
  mindset
- |
  mineable
- |
  minefield
- |
  minelayer
- |
  miner
- |
  mineral
- |
  mineralize
- |
  mineralogist
- |
  mineralogy
- |
  Minerva
- |
  minestrone
- |
  minesweeper
- |
  mingily
- |
  mingle
- |
  mingler
- |
  mingy
- |
  miniature
- |
  miniaturist
- |
  miniaturize
- |
  minibike
- |
  minibus
- |
  minicam
- |
  minicomputer
- |
  minim
- |
  minima
- |
  minimal
- |
  minimalism
- |
  minimalist
- |
  minimally
- |
  minimise
- |
  minimization
- |
  minimize
- |
  minimizer
- |
  minimum
- |
  mining
- |
  minion
- |
  miniscule
- |
  miniseries
- |
  miniskirt
- |
  miniskirted
- |
  minister
- |
  ministerial
- |
  ministrant
- |
  ministration
- |
  ministrative
- |
  ministry
- |
  minivan
- |
  Minneapolis
- |
  minnesinger
- |
  Minnesota
- |
  Minnesotan
- |
  Minnie
- |
  minnow
- |
  Minoan
- |
  minor
- |
  Minorca
- |
  Minorcan
- |
  minority
- |
  minors
- |
  Minotaur
- |
  minoxidil
- |
  Minsk
- |
  minster
- |
  minstrel
- |
  minstrelsy
- |
  mintage
- |
  minter
- |
  minting
- |
  minty
- |
  minuend
- |
  minuet
- |
  Minuit
- |
  minus
- |
  minuscular
- |
  minuscule
- |
  minute
- |
  minutely
- |
  Minuteman
- |
  minuteman
- |
  minuteness
- |
  minutes
- |
  minutia
- |
  minutiae
- |
  minxish
- |
  minyan
- |
  minyanim
- |
  Miocene
- |
  Mirach
- |
  miracle
- |
  miraculous
- |
  miraculously
- |
  mirage
- |
  Miranda
- |
  Mirfak
- |
  Miriam
- |
  mirin
- |
  mirror
- |
  mirrored
- |
  mirth
- |
  mirthful
- |
  mirthfully
- |
  mirthfulness
- |
  mirthless
- |
  mirthlessly
- |
  misaddress
- |
  misadventure
- |
  misadvise
- |
  misaligned
- |
  misalignment
- |
  misalliance
- |
  misallocate
- |
  misally
- |
  misanthrope
- |
  misanthropic
- |
  misanthropy
- |
  misapply
- |
  misapprehend
- |
  misattribute
- |
  misbegotten
- |
  misbehave
- |
  misbehaver
- |
  misbehavior
- |
  misbelieve
- |
  misbeliever
- |
  misbrand
- |
  miscalculate
- |
  miscall
- |
  miscarriage
- |
  miscarry
- |
  miscast
- |
  miscellany
- |
  mischance
- |
  mischief
- |
  mischievous
- |
  miscibility
- |
  miscible
- |
  misclassify
- |
  misconceive
- |
  misconceiver
- |
  misconduct
- |
  misconstrue
- |
  miscopy
- |
  miscount
- |
  miscreant
- |
  miscue
- |
  misdate
- |
  misdeal
- |
  misdealt
- |
  misdeed
- |
  misdefine
- |
  misdemeanor
- |
  misdemeanour
- |
  misdiagnose
- |
  misdiagnosis
- |
  misdial
- |
  misdid
- |
  misdirect
- |
  misdirection
- |
  misdo
- |
  misdoer
- |
  misdoing
- |
  misdone
- |
  miseducate
- |
  misemploy
- |
  miser
- |
  miserable
- |
  miserably
- |
  miserliness
- |
  miserly
- |
  misery
- |
  misestimate
- |
  misfeasance
- |
  misfile
- |
  misfire
- |
  misfit
- |
  misfortune
- |
  misgiving
- |
  misgivings
- |
  misgovern
- |
  misguidance
- |
  misguide
- |
  misguided
- |
  misguidedly
- |
  mishandle
- |
  mishap
- |
  mishear
- |
  misheard
- |
  mishmash
- |
  misidentify
- |
  misinform
- |
  misinterpret
- |
  misjudge
- |
  misjudgment
- |
  Miskito
- |
  mislabel
- |
  mislaid
- |
  mislay
- |
  mislead
- |
  misleading
- |
  misleadingly
- |
  misled
- |
  mislike
- |
  mismanage
- |
  mismatch
- |
  mismatched
- |
  mismate
- |
  misname
- |
  misnomer
- |
  misnumber
- |
  misogamist
- |
  misogamy
- |
  misogynist
- |
  misogynistic
- |
  misogynous
- |
  misogyny
- |
  misorient
- |
  misperceive
- |
  misplace
- |
  misplaced
- |
  misplacement
- |
  misplay
- |
  misprint
- |
  misprision
- |
  mispronounce
- |
  misquotation
- |
  misquote
- |
  misread
- |
  misreading
- |
  misreckon
- |
  misregister
- |
  misremember
- |
  misreport
- |
  misrepresent
- |
  misrule
- |
  missal
- |
  missend
- |
  misshape
- |
  misshapen
- |
  misshapenly
- |
  missile
- |
  missilery
- |
  missilry
- |
  missing
- |
  mission
- |
  missionary
- |
  missioner
- |
  missis
- |
  Mississauga
- |
  Mississippi
- |
  missive
- |
  Missouri
- |
  Missourian
- |
  misspeak
- |
  misspell
- |
  misspelling
- |
  misspelt
- |
  misspend
- |
  misspent
- |
  misstate
- |
  misstatement
- |
  misstep
- |
  missus
- |
  mistakable
- |
  mistake
- |
  mistaken
- |
  mistakenly
- |
  mistaker
- |
  Mister
- |
  mister
- |
  misthrew
- |
  misthrow
- |
  misthrown
- |
  mistily
- |
  mistime
- |
  mistiness
- |
  mistitle
- |
  mistletoe
- |
  mistook
- |
  mistral
- |
  mistranslate
- |
  mistreat
- |
  mistreatment
- |
  Mistress
- |
  mistress
- |
  mistrial
- |
  mistrust
- |
  mistrustful
- |
  misty
- |
  mistype
- |
  misusage
- |
  misuse
- |
  misvalue
- |
  misword
- |
  miswrite
- |
  Mitchell
- |
  miter
- |
  Mitford
- |
  Mithridates
- |
  mitigable
- |
  mitigate
- |
  mitigating
- |
  mitigation
- |
  mitigative
- |
  mitigator
- |
  mitigatory
- |
  mitochondria
- |
  mitoses
- |
  mitosis
- |
  mitotic
- |
  mitotically
- |
  mitre
- |
  mitten
- |
  Mitterrand
- |
  Mitty
- |
  Mitzi
- |
  mitzvah
- |
  mitzvoth
- |
  mixable
- |
  mixed
- |
  mixer
- |
  mixing
- |
  mixologist
- |
  mixology
- |
  Mixtec
- |
  mixture
- |
  mixup
- |
  Mizar
- |
  mizen
- |
  mizenmast
- |
  mizzen
- |
  mizzenmast
- |
  mizzensail
- |
  mnemonic
- |
  mnemonically
- |
  Moabite
- |
  moaner
- |
  Mobile
- |
  mobile
- |
  mobilise
- |
  mobility
- |
  mobilization
- |
  mobilize
- |
  mobilizer
- |
  mobster
- |
  moccasin
- |
  mocha
- |
  mocker
- |
  mockery
- |
  mocking
- |
  mockingbird
- |
  mockingly
- |
  mockup
- |
  modal
- |
  modality
- |
  modally
- |
  model
- |
  modeler
- |
  modeling
- |
  modelling
- |
  modem
- |
  Modena
- |
  moderate
- |
  moderately
- |
  moderateness
- |
  moderation
- |
  moderator
- |
  modern
- |
  moderne
- |
  modernise
- |
  Modernism
- |
  modernism
- |
  modernist
- |
  modernistic
- |
  modernity
- |
  modernize
- |
  modernizer
- |
  modernizing
- |
  modernly
- |
  modernness
- |
  modest
- |
  modestly
- |
  Modesto
- |
  modesty
- |
  modicum
- |
  modification
- |
  modifier
- |
  modify
- |
  Modigliani
- |
  modish
- |
  modishly
- |
  modishness
- |
  modiste
- |
  modular
- |
  modularized
- |
  modulate
- |
  modulation
- |
  modulator
- |
  modulatory
- |
  module
- |
  Mogadiscio
- |
  Mogadishu
- |
  Moghul
- |
  Mogilyov
- |
  Mogul
- |
  mogul
- |
  mohair
- |
  Mohammed
- |
  Mohammedan
- |
  Mohave
- |
  Mohawk
- |
  Mohegan
- |
  Mohican
- |
  moiety
- |
  moiler
- |
  moire
- |
  moist
- |
  moisten
- |
  moistener
- |
  moistly
- |
  moistness
- |
  moisture
- |
  moisturiser
- |
  moisturize
- |
  moisturizer
- |
  Mojave
- |
  molal
- |
  molality
- |
  molar
- |
  molasses
- |
  moldable
- |
  Moldavia
- |
  Moldavian
- |
  moldboard
- |
  molder
- |
  moldering
- |
  moldiness
- |
  molding
- |
  Moldova
- |
  Moldovan
- |
  moldy
- |
  molecular
- |
  molecularity
- |
  molecule
- |
  molehill
- |
  moleskin
- |
  molest
- |
  molestation
- |
  molester
- |
  Moliere
- |
  Mollie
- |
  mollie
- |
  mollifier
- |
  mollify
- |
  mollusc
- |
  molluscan
- |
  mollusk
- |
  molluskan
- |
  Molly
- |
  molly
- |
  mollycoddle
- |
  mollycoddler
- |
  Molnar
- |
  Molokai
- |
  molten
- |
  molter
- |
  Molucca
- |
  Moluccan
- |
  Moluccas
- |
  molybdenum
- |
  Mombasa
- |
  moment
- |
  momenta
- |
  momentarily
- |
  momentary
- |
  momentous
- |
  momentously
- |
  momentum
- |
  momma
- |
  Mommsen
- |
  mommy
- |
  Monacan
- |
  Monaco
- |
  monad
- |
  monadic
- |
  monadism
- |
  monadnock
- |
  monarch
- |
  monarchal
- |
  monarchial
- |
  monarchic
- |
  monarchical
- |
  monarchism
- |
  monarchist
- |
  monarchistic
- |
  monarchy
- |
  monasterial
- |
  monastery
- |
  monastic
- |
  monastical
- |
  monastically
- |
  monasticism
- |
  monaural
- |
  monaurally
- |
  Mondale
- |
  Monday
- |
  Mondrian
- |
  Monegasque
- |
  Monet
- |
  monetarily
- |
  monetarism
- |
  monetarist
- |
  monetaristic
- |
  monetary
- |
  monetization
- |
  monetize
- |
  money
- |
  moneybag
- |
  moneybags
- |
  moneyed
- |
  moneylender
- |
  moneymaker
- |
  moneymaking
- |
  moneys
- |
  mongeese
- |
  monger
- |
  mongo
- |
  Mongol
- |
  Mongolia
- |
  Mongolian
- |
  Mongolic
- |
  Mongolism
- |
  mongolism
- |
  Mongoloid
- |
  mongoloid
- |
  mongoose
- |
  mongrel
- |
  Monica
- |
  monicker
- |
  monied
- |
  monies
- |
  moniker
- |
  monikered
- |
  monism
- |
  monist
- |
  monistic
- |
  monition
- |
  monitor
- |
  monitory
- |
  monkey
- |
  monkeyshine
- |
  monkeyshines
- |
  monkish
- |
  monkishly
- |
  monkshood
- |
  Monmouth
- |
  Monoceros
- |
  monochrome
- |
  monochromic
- |
  monocle
- |
  monocled
- |
  monoclinal
- |
  monocline
- |
  monoclonal
- |
  monocoque
- |
  monocot
- |
  monocular
- |
  monocultural
- |
  monoculture
- |
  monodic
- |
  monodical
- |
  monodist
- |
  monody
- |
  monofilament
- |
  monogamist
- |
  monogamous
- |
  monogamously
- |
  monogamy
- |
  monogram
- |
  monogrammed
- |
  monograph
- |
  monographer
- |
  monographic
- |
  monographist
- |
  monolingual
- |
  monolith
- |
  monolithic
- |
  monolog
- |
  monologist
- |
  monologue
- |
  monologuist
- |
  monomania
- |
  monomaniac
- |
  monomaniacal
- |
  monomer
- |
  monomeric
- |
  monomial
- |
  Monongahela
- |
  monophonic
- |
  monoplane
- |
  monopolise
- |
  monopolist
- |
  monopolistic
- |
  monopolize
- |
  monopolizer
- |
  Monopoly
- |
  monopoly
- |
  monorail
- |
  monosyllabic
- |
  monosyllable
- |
  monotheism
- |
  monotheist
- |
  monotheistic
- |
  monotone
- |
  monotonous
- |
  monotonously
- |
  monotony
- |
  monotype
- |
  monotypic
- |
  monovalence
- |
  monovalency
- |
  monovalent
- |
  monoxide
- |
  monozygotic
- |
  Monroe
- |
  Monrovia
- |
  monseigneur
- |
  Monsieur
- |
  monsieur
- |
  Monsignor
- |
  monsignor
- |
  monsignori
- |
  monsoon
- |
  monsoonal
- |
  monster
- |
  monstrance
- |
  monstrosity
- |
  monstrous
- |
  monstrously
- |
  montage
- |
  Montagnais
- |
  Montaigne
- |
  Montana
- |
  Montanan
- |
  Montcalm
- |
  Monte
- |
  Montenegran
- |
  Montenegrin
- |
  Montenegro
- |
  Monterey
- |
  Monterrey
- |
  Montesquieu
- |
  Montessori
- |
  Monteverdi
- |
  Montevideo
- |
  Montezuma
- |
  Montgomery
- |
  month
- |
  monthlong
- |
  monthly
- |
  Monticello
- |
  Montpelier
- |
  Montreal
- |
  Montserrat
- |
  Monty
- |
  monument
- |
  monumental
- |
  monumentally
- |
  mooch
- |
  moocher
- |
  moodily
- |
  moodiness
- |
  moody
- |
  moonbeam
- |
  moonless
- |
  moonlight
- |
  moonlighter
- |
  moonlighting
- |
  moonlit
- |
  moonscape
- |
  moonshine
- |
  moonshiner
- |
  moonshot
- |
  moonstone
- |
  moonstruck
- |
  moonwalk
- |
  moony
- |
  moorage
- |
  Moore
- |
  mooring
- |
  moorings
- |
  Moorish
- |
  moorland
- |
  moose
- |
  moped
- |
  moper
- |
  mopey
- |
  mopish
- |
  mopishly
- |
  mopper
- |
  moppet
- |
  moraine
- |
  moral
- |
  morale
- |
  moralist
- |
  moralistic
- |
  morality
- |
  moralization
- |
  moralize
- |
  moralizer
- |
  moralizing
- |
  moralizingly
- |
  morally
- |
  morals
- |
  morass
- |
  moratoria
- |
  moratorium
- |
  Moravia
- |
  Moravian
- |
  moray
- |
  morbid
- |
  morbidity
- |
  morbidly
- |
  morbidness
- |
  mordacious
- |
  mordaciously
- |
  mordacity
- |
  mordancy
- |
  mordant
- |
  mordantly
- |
  Mordecai
- |
  mordent
- |
  Morea
- |
  Morean
- |
  morel
- |
  Morelia
- |
  Morelos
- |
  moreover
- |
  mores
- |
  Morgan
- |
  morgue
- |
  moribund
- |
  moribundity
- |
  moribundly
- |
  Morison
- |
  Morisot
- |
  Mormon
- |
  Mormonism
- |
  morning
- |
  Moroccan
- |
  Morocco
- |
  morocco
- |
  Moron
- |
  moron
- |
  Moroni
- |
  moronic
- |
  moronically
- |
  morose
- |
  morosely
- |
  moroseness
- |
  morph
- |
  morpheme
- |
  morphemic
- |
  Morpheus
- |
  morphia
- |
  morphine
- |
  morphing
- |
  morphogenic
- |
  morphologic
- |
  morphologist
- |
  morphology
- |
  Morris
- |
  morris
- |
  Morrison
- |
  morrow
- |
  Morse
- |
  morsel
- |
  mortal
- |
  mortality
- |
  mortally
- |
  mortar
- |
  mortarboard
- |
  mortgage
- |
  mortgageable
- |
  mortgagee
- |
  mortgager
- |
  mortgagor
- |
  mortice
- |
  mortician
- |
  mortify
- |
  mortifying
- |
  mortifyingly
- |
  Mortimer
- |
  mortise
- |
  mortiser
- |
  mortmain
- |
  Morton
- |
  mortuary
- |
  Mosaic
- |
  mosaic
- |
  mosaicist
- |
  mosaicked
- |
  Moscow
- |
  Mosel
- |
  Moselle
- |
  Moses
- |
  mosey
- |
  Moslem
- |
  mosque
- |
  Mosquito
- |
  mosquito
- |
  mossback
- |
  mossbacked
- |
  mossiness
- |
  mossy
- |
  mostly
- |
  Mosul
- |
  motel
- |
  motet
- |
  mothball
- |
  mothballs
- |
  mother
- |
  motherboard
- |
  motherfucker
- |
  motherhood
- |
  mothering
- |
  Motherland
- |
  motherland
- |
  motherless
- |
  motherliness
- |
  motherly
- |
  mothproof
- |
  motif
- |
  motile
- |
  motility
- |
  motion
- |
  motionless
- |
  motionlessly
- |
  motivate
- |
  motivated
- |
  motivation
- |
  motivational
- |
  motivator
- |
  motive
- |
  motiveless
- |
  motley
- |
  motocross
- |
  motor
- |
  motorbike
- |
  motorboat
- |
  motorcade
- |
  motorcar
- |
  motorcycle
- |
  motorcyclist
- |
  motoring
- |
  motorist
- |
  motorization
- |
  motorize
- |
  motorized
- |
  motorman
- |
  motormouth
- |
  motortruck
- |
  motorway
- |
  mottle
- |
  mottled
- |
  mottling
- |
  motto
- |
  mould
- |
  moulder
- |
  moulding
- |
  mouldy
- |
  Moulmein
- |
  moult
- |
  mound
- |
  Mount
- |
  mount
- |
  mountable
- |
  mountain
- |
  mountaineer
- |
  mountainous
- |
  mountainside
- |
  mountaintop
- |
  mountainy
- |
  Mountbatten
- |
  mountebank
- |
  mounted
- |
  mounter
- |
  Mountie
- |
  mounting
- |
  Mounty
- |
  mourn
- |
  Mourne
- |
  mourner
- |
  mournful
- |
  mournfully
- |
  mournfulness
- |
  mourning
- |
  mouse
- |
  mousepad
- |
  mouser
- |
  mousetrap
- |
  mousey
- |
  mousiness
- |
  moussaka
- |
  mousse
- |
  Moussorgsky
- |
  moustache
- |
  moustached
- |
  mousy
- |
  mouth
- |
  mouthed
- |
  mouthful
- |
  mouthiness
- |
  mouthpart
- |
  mouthpiece
- |
  mouthwash
- |
  mouthy
- |
  mouton
- |
  movability
- |
  movable
- |
  movableness
- |
  movables
- |
  movably
- |
  moveable
- |
  moved
- |
  movement
- |
  mover
- |
  movie
- |
  moviedom
- |
  movies
- |
  moving
- |
  movingly
- |
  mower
- |
  moxie
- |
  Moyle
- |
  Mozambican
- |
  Mozambique
- |
  Mozart
- |
  mozzarella
- |
  Mubarak
- |
  mucilage
- |
  mucilaginous
- |
  muckrake
- |
  muckraker
- |
  muckraking
- |
  mucky
- |
  mucosa
- |
  mucosae
- |
  mucosity
- |
  mucous
- |
  mucus
- |
  muddied
- |
  muddily
- |
  muddiness
- |
  muddle
- |
  muddled
- |
  muddleheaded
- |
  muddler
- |
  muddy
- |
  mudflat
- |
  mudguard
- |
  mudroom
- |
  mudslide
- |
  mudslinger
- |
  mudslinging
- |
  Muenster
- |
  muenster
- |
  muesli
- |
  muezzin
- |
  muffin
- |
  muffle
- |
  muffled
- |
  muffler
- |
  mufti
- |
  Mugabe
- |
  mugful
- |
  mugger
- |
  mugginess
- |
  mugging
- |
  muggy
- |
  Mughal
- |
  mugshot
- |
  mugwump
- |
  mugwumpery
- |
  Muhammad
- |
  Muhammadan
- |
  Muharram
- |
  mujahedeen
- |
  mujahedin
- |
  mujahideen
- |
  mujahidin
- |
  Mukden
- |
  mukluk
- |
  mulatto
- |
  mulberry
- |
  mulch
- |
  mulct
- |
  muleskinner
- |
  muleteer
- |
  muliebrity
- |
  mulish
- |
  mulishly
- |
  mulishness
- |
  mulla
- |
  mullah
- |
  mullein
- |
  mullen
- |
  mullet
- |
  mulligan
- |
  mulligatawny
- |
  mullion
- |
  mullioned
- |
  Mulroney
- |
  Multan
- |
  multicolor
- |
  multicolored
- |
  multiethnic
- |
  multifaceted
- |
  multifamily
- |
  multifarious
- |
  multiform
- |
  multiformity
- |
  multilane
- |
  multilateral
- |
  multilayered
- |
  multilevel
- |
  multilingual
- |
  multimedia
- |
  multiparous
- |
  multiple
- |
  multiplex
- |
  multiplexer
- |
  multiplexity
- |
  multiplexor
- |
  multiplicand
- |
  multiplicity
- |
  multiplier
- |
  multiply
- |
  multipurpose
- |
  multiracial
- |
  multisense
- |
  multistage
- |
  multistory
- |
  multitask
- |
  multitasking
- |
  multitude
- |
  multiunit
- |
  multiuse
- |
  multivalence
- |
  multivalency
- |
  multivalent
- |
  multivitamin
- |
  Mumbai
- |
  mumble
- |
  mumbler
- |
  mumbletypeg
- |
  mumbly
- |
  mummer
- |
  mummery
- |
  mummify
- |
  mummy
- |
  mumps
- |
  munch
- |
  munchies
- |
  mundane
- |
  mundanely
- |
  mundaneness
- |
  mundanity
- |
  Munich
- |
  municipal
- |
  municipality
- |
  municipalize
- |
  municipally
- |
  munificence
- |
  munificent
- |
  munificently
- |
  muniment
- |
  muniments
- |
  munition
- |
  munitioner
- |
  munitions
- |
  Munro
- |
  Munster
- |
  mural
- |
  muralist
- |
  Murat
- |
  Murcia
- |
  Murcian
- |
  murder
- |
  murderer
- |
  murderess
- |
  murderous
- |
  murderously
- |
  Murdoch
- |
  murex
- |
  murices
- |
  Muriel
- |
  murkily
- |
  murkiness
- |
  murky
- |
  Murmansk
- |
  murmur
- |
  murmurer
- |
  murmuring
- |
  murmurous
- |
  murrain
- |
  Murray
- |
  Murrow
- |
  Murrumbidgee
- |
  Musca
- |
  Muscat
- |
  muscat
- |
  muscatel
- |
  muscle
- |
  musclebound
- |
  muscled
- |
  Muscovite
- |
  Muscovy
- |
  muscular
- |
  muscularity
- |
  muscularly
- |
  musculature
- |
  muser
- |
  Muses
- |
  musette
- |
  museum
- |
  mushiness
- |
  mushroom
- |
  mushrooming
- |
  mushy
- |
  music
- |
  musical
- |
  musicale
- |
  musicality
- |
  musically
- |
  musician
- |
  musicianly
- |
  musicianship
- |
  musicologist
- |
  musicology
- |
  musing
- |
  musingly
- |
  muskeg
- |
  muskellunge
- |
  musket
- |
  musketeer
- |
  musketry
- |
  muskie
- |
  muskiness
- |
  muskmelon
- |
  Muskogean
- |
  Muskogee
- |
  muskox
- |
  muskoxen
- |
  muskrat
- |
  musky
- |
  Muslim
- |
  muslin
- |
  mussel
- |
  mussily
- |
  mussiness
- |
  Mussolini
- |
  Mussorgsky
- |
  mussy
- |
  mustache
- |
  mustached
- |
  mustachio
- |
  mustang
- |
  mustard
- |
  mustardy
- |
  muster
- |
  musth
- |
  mustily
- |
  mustiness
- |
  musty
- |
  mutability
- |
  mutable
- |
  mutableness
- |
  mutably
- |
  mutagen
- |
  mutagenesis
- |
  mutagenic
- |
  mutant
- |
  mutate
- |
  mutation
- |
  mutational
- |
  mutationally
- |
  mutative
- |
  muted
- |
  mutely
- |
  muteness
- |
  mutilate
- |
  mutilated
- |
  mutilation
- |
  mutilative
- |
  mutilator
- |
  mutineer
- |
  mutinous
- |
  mutinously
- |
  mutiny
- |
  mutism
- |
  mutter
- |
  mutterer
- |
  mutton
- |
  muttonchops
- |
  muttony
- |
  mutual
- |
  mutualism
- |
  mutualist
- |
  mutualistic
- |
  mutuality
- |
  mutually
- |
  muumuu
- |
  Muzak
- |
  muzzily
- |
  muzziness
- |
  muzzle
- |
  muzzleloader
- |
  muzzy
- |
  Mwanza
- |
  myalgia
- |
  myalgic
- |
  Myanma
- |
  Myanmar
- |
  myasthenia
- |
  myasthenic
- |
  mycelia
- |
  mycelial
- |
  mycelium
- |
  Mycenae
- |
  Mycenaean
- |
  mycological
- |
  mycologist
- |
  mycology
- |
  myelin
- |
  myeline
- |
  myelitis
- |
  myeloma
- |
  myelomata
- |
  Mykolayiv
- |
  Mylar
- |
  Myles
- |
  mynah
- |
  myocardia
- |
  myocardial
- |
  myocardium
- |
  myological
- |
  myologist
- |
  myology
- |
  myopia
- |
  myopic
- |
  myopically
- |
  myosin
- |
  myriad
- |
  myriapod
- |
  myrmidon
- |
  Myrna
- |
  Myron
- |
  myrrh
- |
  Myrtle
- |
  myrtle
- |
  myself
- |
  Mysore
- |
  mystagogical
- |
  mystagogue
- |
  mystagogy
- |
  mysteries
- |
  mysterious
- |
  mysteriously
- |
  mystery
- |
  mystic
- |
  mystical
- |
  mystically
- |
  mysticalness
- |
  mysticism
- |
  mystify
- |
  mystifying
- |
  mystifyingly
- |
  mystique
- |
  mythic
- |
  mythical
- |
  mythically
- |
  mythicism
- |
  mythicist
- |
  mythicize
- |
  mythmaker
- |
  mythmaking
- |
  mythologer
- |
  mythologic
- |
  mythological
- |
  mythologist
- |
  mythologize
- |
  mythology
- |
  mythomane
- |
  mythomania
- |
  mythomaniac
- |
  Myukolayiv
- |
  Nabataea
- |
  Nabataean
- |
  Nabatea
- |
  Nabatean
- |
  nabob
- |
  Nabokov
- |
  nacelle
- |
  nacho
- |
  nacre
- |
  nacreous
- |
  NaDene
- |
  Nader
- |
  Nadia
- |
  Nadine
- |
  nadir
- |
  naevi
- |
  naevus
- |
  Nagasaki
- |
  nagger
- |
  nagging
- |
  naggingly
- |
  Nagoya
- |
  Nagpur
- |
  Nahuatl
- |
  Nahum
- |
  Naiad
- |
  naiad
- |
  naiades
- |
  nailbrush
- |
  nailer
- |
  nainsook
- |
  Naipaul
- |
  naira
- |
  Nairobi
- |
  naive
- |
  naively
- |
  naiveness
- |
  naivete
- |
  naivety
- |
  naked
- |
  nakedly
- |
  nakedness
- |
  nakfa
- |
  namable
- |
  nameable
- |
  namedrop
- |
  namedropping
- |
  nameless
- |
  namelessly
- |
  namelessness
- |
  namely
- |
  nameplate
- |
  namer
- |
  namesake
- |
  Namibia
- |
  Namibian
- |
  Nampula
- |
  Nanchang
- |
  Nancy
- |
  Nanette
- |
  Nanjing
- |
  nankeen
- |
  nankin
- |
  Nanking
- |
  Nannette
- |
  nanny
- |
  nanometer
- |
  nanosecond
- |
  nanotube
- |
  Nansen
- |
  Nantes
- |
  Nantucket
- |
  Nantucketer
- |
  Naomi
- |
  napalm
- |
  napery
- |
  naphtha
- |
  naphthalene
- |
  naphthous
- |
  Napier
- |
  napkin
- |
  Naples
- |
  napless
- |
  Napoleon
- |
  napoleon
- |
  Napoleonic
- |
  napped
- |
  napper
- |
  nappy
- |
  Napster
- |
  narcissi
- |
  narcissism
- |
  narcissist
- |
  narcissistic
- |
  Narcissus
- |
  narcissus
- |
  narcolepsy
- |
  narcoleptic
- |
  narcoses
- |
  narcosis
- |
  narcotic
- |
  narcotically
- |
  narcotism
- |
  narcotize
- |
  nares
- |
  naris
- |
  Narraganset
- |
  Narragansett
- |
  narrate
- |
  narration
- |
  narrative
- |
  narrator
- |
  narrow
- |
  narrowly
- |
  narrowness
- |
  narrows
- |
  narthex
- |
  narwhal
- |
  nasal
- |
  nasality
- |
  nasalization
- |
  nasalize
- |
  nasally
- |
  nascence
- |
  nascency
- |
  nascent
- |
  Nashik
- |
  Nashua
- |
  Nashville
- |
  Nasik
- |
  Nassau
- |
  Nasser
- |
  nastily
- |
  nastiness
- |
  nasturtium
- |
  nasty
- |
  Natal
- |
  natal
- |
  Natalie
- |
  natality
- |
  natatorium
- |
  Natchez
- |
  nates
- |
  Nathan
- |
  Nathanael
- |
  Nathaniel
- |
  Natick
- |
  Nation
- |
  nation
- |
  national
- |
  nationalise
- |
  nationalism
- |
  nationalist
- |
  nationality
- |
  nationalize
- |
  nationalized
- |
  nationalizer
- |
  nationally
- |
  nationhood
- |
  nationwide
- |
  native
- |
  nativism
- |
  nativist
- |
  nativistic
- |
  Nativity
- |
  nativity
- |
  natter
- |
  natterer
- |
  nattily
- |
  nattiness
- |
  natty
- |
  natural
- |
  naturalism
- |
  naturalist
- |
  naturalistic
- |
  naturalize
- |
  naturalized
- |
  naturally
- |
  naturalness
- |
  nature
- |
  natured
- |
  naturism
- |
  naturist
- |
  naturopath
- |
  naturopathic
- |
  naturopathy
- |
  Naugahyde
- |
  naught
- |
  naughtily
- |
  naughtiness
- |
  naughty
- |
  Nauru
- |
  Nauruan
- |
  nausea
- |
  nauseate
- |
  nauseated
- |
  nauseating
- |
  nauseatingly
- |
  nauseation
- |
  nauseous
- |
  nauseously
- |
  nauseousness
- |
  nautical
- |
  nautically
- |
  nautili
- |
  nautilus
- |
  Navaho
- |
  Navajo
- |
  naval
- |
  Navarre
- |
  navel
- |
  navigability
- |
  navigable
- |
  navigate
- |
  navigation
- |
  navigational
- |
  navigator
- |
  Navratilova
- |
  Nayarit
- |
  naysayer
- |
  Nazarene
- |
  Nazareth
- |
  Naziism
- |
  Nazism
- |
  Ndola
- |
  Neanderthal
- |
  neanderthal
- |
  Neapolis
- |
  Neapolitan
- |
  nearby
- |
  nearish
- |
  nearly
- |
  nearness
- |
  nearsighted
- |
  neaten
- |
  neath
- |
  neatly
- |
  neatness
- |
  nebbich
- |
  nebbish
- |
  Nebraska
- |
  Nebraskan
- |
  nebula
- |
  nebulae
- |
  nebular
- |
  nebulization
- |
  nebulize
- |
  nebulizer
- |
  nebulosity
- |
  nebulous
- |
  nebulously
- |
  nebulousness
- |
  necessarily
- |
  necessary
- |
  necessitate
- |
  necessitous
- |
  necessity
- |
  necked
- |
  neckerchief
- |
  necking
- |
  necklace
- |
  necklacing
- |
  neckline
- |
  necktie
- |
  neckwear
- |
  necrologic
- |
  necrological
- |
  necrologist
- |
  necrology
- |
  necromancer
- |
  necromancy
- |
  necromantic
- |
  necrophile
- |
  necrophilia
- |
  necrophiliac
- |
  necrophilic
- |
  necrophilism
- |
  necrophilist
- |
  necropoleis
- |
  necropoles
- |
  necropoli
- |
  necropolis
- |
  necroses
- |
  necrosis
- |
  necrotic
- |
  nectar
- |
  nectarine
- |
  nectarous
- |
  needful
- |
  needfully
- |
  needfulness
- |
  neediness
- |
  needle
- |
  needlepoint
- |
  needler
- |
  needless
- |
  needlessly
- |
  needlessness
- |
  needlewoman
- |
  needlework
- |
  needs
- |
  needy
- |
  nefarious
- |
  nefariously
- |
  Nefertiti
- |
  negate
- |
  negation
- |
  negative
- |
  negatively
- |
  negativeness
- |
  negativism
- |
  negativist
- |
  negativistic
- |
  negativity
- |
  negatory
- |
  negatron
- |
  Negev
- |
  neglect
- |
  neglected
- |
  neglecter
- |
  neglectful
- |
  neglectfully
- |
  neglige
- |
  negligee
- |
  negligence
- |
  negligent
- |
  negligently
- |
  negligible
- |
  negligibly
- |
  negotiable
- |
  negotiant
- |
  negotiate
- |
  negotiation
- |
  negotiator
- |
  Negress
- |
  Negritude
- |
  negritude
- |
  Negro
- |
  Negroid
- |
  Negros
- |
  Nehemiah
- |
  Nehru
- |
  neigh
- |
  neighbor
- |
  neighborhood
- |
  neighboring
- |
  neighborly
- |
  neighbour
- |
  neighbouring
- |
  neither
- |
  Nellie
- |
  Nelson
- |
  nelson
- |
  nematode
- |
  Nemea
- |
  Nemean
- |
  nemeses
- |
  Nemesis
- |
  nemesis
- |
  neoclassic
- |
  neoclassical
- |
  neocolonial
- |
  neodymium
- |
  neoliberal
- |
  Neolithic
- |
  neolithic
- |
  neological
- |
  neologism
- |
  neologist
- |
  neologize
- |
  neonatal
- |
  neonatally
- |
  neonate
- |
  neonatology
- |
  neophyte
- |
  neoplasm
- |
  neoplastic
- |
  neoprene
- |
  neoteric
- |
  Nepal
- |
  Nepalese
- |
  Nepali
- |
  nepenthe
- |
  nephew
- |
  nephrite
- |
  nephritic
- |
  nephritides
- |
  nephritis
- |
  nephrosis
- |
  nepotism
- |
  nepotist
- |
  nepotistic
- |
  Neptune
- |
  Neptunian
- |
  neptunium
- |
  nerdy
- |
  Nereid
- |
  nereid
- |
  Neronian
- |
  Neruda
- |
  nerve
- |
  nerved
- |
  nerveless
- |
  nervelessly
- |
  nerveracking
- |
  nerves
- |
  nervily
- |
  nerviness
- |
  nervous
- |
  nervously
- |
  nervousness
- |
  nervy
- |
  nescience
- |
  nescient
- |
  nestle
- |
  nestler
- |
  nestling
- |
  Nestor
- |
  nether
- |
  Netherland
- |
  Netherlander
- |
  Netherlands
- |
  nethermost
- |
  netherworld
- |
  netiquette
- |
  Nettie
- |
  netting
- |
  nettle
- |
  nettlesome
- |
  network
- |
  networking
- |
  neural
- |
  neuralgia
- |
  neuralgic
- |
  neurally
- |
  neurasthenia
- |
  neurasthenic
- |
  neuritic
- |
  neuritides
- |
  neuritis
- |
  neurologic
- |
  neurological
- |
  neurologist
- |
  neurology
- |
  neuron
- |
  neuronal
- |
  neurone
- |
  neuronic
- |
  neuroscience
- |
  neuroses
- |
  neurosis
- |
  neurosurgeon
- |
  neurosurgery
- |
  neurotic
- |
  neurotically
- |
  neuter
- |
  neutered
- |
  neutral
- |
  neutralise
- |
  neutralism
- |
  neutralist
- |
  neutrality
- |
  neutralize
- |
  neutralizer
- |
  neutrally
- |
  neutrino
- |
  neutron
- |
  Nevada
- |
  Nevadan
- |
  Nevadian
- |
  Nevelson
- |
  never
- |
  nevermore
- |
  nevertheless
- |
  Nevil
- |
  Neville
- |
  Nevin
- |
  Nevis
- |
  nevus
- |
  Newark
- |
  newbie
- |
  newborn
- |
  Newcastle
- |
  newcomer
- |
  newel
- |
  Newell
- |
  newfangled
- |
  newfound
- |
  Newfoundland
- |
  Newham
- |
  newish
- |
  newly
- |
  newlywed
- |
  newlyweds
- |
  Newman
- |
  newness
- |
  Newport
- |
  Newry
- |
  newsagent
- |
  newsboy
- |
  newscast
- |
  newscaster
- |
  newsdealer
- |
  newsgroup
- |
  newsletter
- |
  newsmagazine
- |
  newsman
- |
  newspaper
- |
  newspaperman
- |
  newspeak
- |
  newsprint
- |
  newsreel
- |
  newsroom
- |
  newsstand
- |
  newsweekly
- |
  newswoman
- |
  newsworthy
- |
  newsy
- |
  Newton
- |
  newton
- |
  Newtonian
- |
  Newtownabbey
- |
  Newtownards
- |
  nextdoor
- |
  nexus
- |
  ngultrum
- |
  ngwee
- |
  niacin
- |
  Niagara
- |
  Niamey
- |
  nibble
- |
  nibbler
- |
  Nicaea
- |
  Nicaean
- |
  Nicaragua
- |
  Nicaraguan
- |
  nicely
- |
  Nicene
- |
  niceness
- |
  niceties
- |
  nicety
- |
  niche
- |
  Nicholas
- |
  nickel
- |
  nickelodeon
- |
  nicker
- |
  Nicklaus
- |
  nickname
- |
  Nicobar
- |
  Nicole
- |
  Nicosia
- |
  nicotine
- |
  nictate
- |
  nictitate
- |
  nictitation
- |
  Niebuhr
- |
  niece
- |
  nielsbohrium
- |
  Nietzsche
- |
  Nietzschean
- |
  nifty
- |
  Niger
- |
  Nigeria
- |
  Nigerian
- |
  Nigerien
- |
  niggard
- |
  niggardly
- |
  nigger
- |
  niggle
- |
  niggler
- |
  niggling
- |
  nigglingly
- |
  night
- |
  nightblind
- |
  nightcap
- |
  nightclothes
- |
  nightclub
- |
  nightdress
- |
  nightfall
- |
  nightgown
- |
  nighthawk
- |
  nightie
- |
  Nightingale
- |
  nightingale
- |
  nightlife
- |
  nightly
- |
  nightmare
- |
  nightmarish
- |
  nights
- |
  nightshade
- |
  nightshirt
- |
  nightspot
- |
  nightstand
- |
  nightstick
- |
  nighttime
- |
  nightwalker
- |
  nightwear
- |
  nighty
- |
  nihilism
- |
  nihilist
- |
  nihilistic
- |
  Nihon
- |
  Niihau
- |
  Nijinsky
- |
  Nikkei
- |
  Niklaus
- |
  Nikolaev
- |
  Nikolayev
- |
  Niles
- |
  Nilgiri
- |
  Nilotic
- |
  Nilsson
- |
  nimbi
- |
  nimble
- |
  nimbleness
- |
  nimbly
- |
  nimbus
- |
  Nimes
- |
  Nimitz
- |
  Nimrod
- |
  nimrod
- |
  nincompoop
- |
  ninefold
- |
  ninepins
- |
  nineteen
- |
  nineteenth
- |
  ninetieth
- |
  ninety
- |
  Nineveh
- |
  ninja
- |
  ninny
- |
  ninth
- |
  Niobe
- |
  niobium
- |
  nipper
- |
  nippers
- |
  nipple
- |
  Nippon
- |
  Nipponese
- |
  nippy
- |
  Nirvana
- |
  nirvana
- |
  Nisan
- |
  Nisei
- |
  nisei
- |
  niter
- |
  nitpick
- |
  nitpicker
- |
  nitpicking
- |
  nitrate
- |
  nitration
- |
  nitre
- |
  nitride
- |
  nitrify
- |
  nitrifying
- |
  nitrite
- |
  nitro
- |
  nitrogen
- |
  nitrogenous
- |
  nitrous
- |
  nitty
- |
  nitwit
- |
  niveous
- |
  Nixon
- |
  Nkrumah
- |
  Nobel
- |
  Nobelist
- |
  nobelium
- |
  nobility
- |
  noble
- |
  nobleman
- |
  nobleness
- |
  noblesse
- |
  noblewoman
- |
  nobly
- |
  nobody
- |
  noctambulism
- |
  noctambulist
- |
  nocturnal
- |
  nocturnally
- |
  nocturne
- |
  nocuous
- |
  nocuously
- |
  nodal
- |
  noddle
- |
  noddy
- |
  nodular
- |
  nodule
- |
  nodus
- |
  noetic
- |
  noggin
- |
  nohow
- |
  noise
- |
  noiseless
- |
  noiselessly
- |
  noisemaker
- |
  noisily
- |
  noisiness
- |
  noisome
- |
  noisomely
- |
  noisomeness
- |
  noisy
- |
  Nolan
- |
  nomad
- |
  nomadic
- |
  nomadically
- |
  nomadism
- |
  nomenclature
- |
  nominal
- |
  nominalism
- |
  nominalist
- |
  nominalistic
- |
  nominally
- |
  nominate
- |
  nomination
- |
  nominative
- |
  nominator
- |
  nominee
- |
  nonabrasive
- |
  nonabsorbent
- |
  nonabusive
- |
  nonacademic
- |
  nonacid
- |
  nonactivated
- |
  nonactive
- |
  nonadaptive
- |
  nonaddicting
- |
  nonaddictive
- |
  nonadherence
- |
  nonadhesive
- |
  nonadjacent
- |
  nonage
- |
  nonagenarian
- |
  nonagon
- |
  nonalcoholic
- |
  nonaligned
- |
  nonalignment
- |
  nonallergic
- |
  nonallied
- |
  nonanalytic
- |
  nonapproved
- |
  nonaromatic
- |
  nonarrival
- |
  nonassertive
- |
  nonathletic
- |
  nonautomatic
- |
  nonbasic
- |
  nonbeliever
- |
  nonbinding
- |
  nonbook
- |
  nonbreakable
- |
  nonburnable
- |
  noncaking
- |
  noncaloric
- |
  noncancerous
- |
  noncandidate
- |
  noncausal
- |
  nonce
- |
  noncellular
- |
  nonchalance
- |
  nonchalant
- |
  nonchalantly
- |
  noncitizen
- |
  nonclerical
- |
  nonclinical
- |
  nonclotting
- |
  noncoherent
- |
  noncoital
- |
  noncom
- |
  noncombat
- |
  noncombatant
- |
  noncommittal
- |
  noncommunist
- |
  noncompeting
- |
  noncompliant
- |
  noncomplying
- |
  nonconductor
- |
  noncorroding
- |
  noncorrosive
- |
  noncredit
- |
  noncriminal
- |
  noncritical
- |
  noncurrent
- |
  noncustodial
- |
  nondairy
- |
  nondeadly
- |
  nondelivery
- |
  nondescript
- |
  nondivisible
- |
  nondogmatic
- |
  nondomestic
- |
  nondominant
- |
  nondramatic
- |
  nondrinker
- |
  nondriver
- |
  nondrug
- |
  nondrying
- |
  nondurable
- |
  noneconomic
- |
  nonedible
- |
  noneffective
- |
  nonelastic
- |
  nonelected
- |
  nonelection
- |
  nonelective
- |
  nonelectric
- |
  noneligible
- |
  nonemergency
- |
  nonemotional
- |
  nonentity
- |
  nones
- |
  nonessential
- |
  nonesuch
- |
  nonetheless
- |
  nonethical
- |
  nonevent
- |
  nonexclusive
- |
  nonexempt
- |
  nonexistence
- |
  nonexistent
- |
  nonexplosive
- |
  nonextinct
- |
  nonfactual
- |
  nonfading
- |
  nonfarm
- |
  nonfascist
- |
  nonfat
- |
  nonfatal
- |
  nonfattening
- |
  nonfeasance
- |
  nonfederated
- |
  nonferrous
- |
  nonfiction
- |
  nonfictional
- |
  nonflammable
- |
  nonflexible
- |
  nonflowering
- |
  nonflying
- |
  nonfood
- |
  nonfreezing
- |
  nongaseous
- |
  nongraded
- |
  nongranular
- |
  nongreasy
- |
  nonhazardous
- |
  nonhero
- |
  nonhuman
- |
  nonidentical
- |
  nonillion
- |
  nonillionth
- |
  noninclusive
- |
  noninductive
- |
  noninfected
- |
  noninflected
- |
  noninvasive
- |
  nonionizing
- |
  nonissue
- |
  nonjoiner
- |
  nonjudicial
- |
  nonkosher
- |
  nonlegal
- |
  nonlethal
- |
  nonlinear
- |
  nonliterary
- |
  nonliving
- |
  nonlogical
- |
  nonmagnetic
- |
  nonmalicious
- |
  nonmalignant
- |
  nonmaterial
- |
  nonmedical
- |
  nonmember
- |
  nonmetal
- |
  nonmetallic
- |
  nonmigratory
- |
  nonmilitant
- |
  nonmilitary
- |
  nonmoral
- |
  nonmotile
- |
  nonmoving
- |
  nonnarcotic
- |
  nonnative
- |
  nonnegative
- |
  nonnuclear
- |
  nonnumerical
- |
  nonobjective
- |
  nonobservant
- |
  nonofficial
- |
  nonoily
- |
  nonoperative
- |
  nonorganic
- |
  nonorthodox
- |
  nonparallel
- |
  nonparasitic
- |
  nonpareil
- |
  nonpartisan
- |
  nonpaternal
- |
  nonpaying
- |
  nonpayment
- |
  nonpermanent
- |
  nonpermeable
- |
  nonperson
- |
  nonphysical
- |
  nonplus
- |
  nonplussed
- |
  nonpoisonous
- |
  nonpolar
- |
  nonpolitical
- |
  nonpolluting
- |
  nonporous
- |
  nonpregnant
- |
  nonprofit
- |
  nonprotein
- |
  nonpublic
- |
  nonracial
- |
  nonrandom
- |
  nonreactive
- |
  nonreader
- |
  nonreceipt
- |
  nonrecurrent
- |
  nonrecurring
- |
  nonreligious
- |
  nonrenewable
- |
  nonresidence
- |
  nonresident
- |
  nonresidual
- |
  nonresistant
- |
  nonrhythmic
- |
  nonrigid
- |
  nonruminant
- |
  nonrural
- |
  nonsalable
- |
  nonsalaried
- |
  nonscheduled
- |
  nonscientist
- |
  nonscoring
- |
  nonseasonal
- |
  nonsectarian
- |
  nonsecular
- |
  nonselective
- |
  nonself
- |
  nonsense
- |
  nonsensical
- |
  nonsensitive
- |
  nonsexist
- |
  nonsexual
- |
  nonsinkable
- |
  nonsked
- |
  nonskid
- |
  nonslip
- |
  nonsmoker
- |
  nonsmoking
- |
  nonsocial
- |
  nonspeaking
- |
  nonspecific
- |
  nonspherical
- |
  nonspiritual
- |
  nonstaining
- |
  nonstandard
- |
  nonstarter
- |
  nonsteroidal
- |
  nonstick
- |
  nonsticking
- |
  nonstop
- |
  nonstrategic
- |
  nonstriking
- |
  nonsuccess
- |
  nonsuch
- |
  nonsuit
- |
  nonsupport
- |
  nonsurgical
- |
  nonswimmer
- |
  nontalkative
- |
  nontaxable
- |
  nonteaching
- |
  nontechnical
- |
  nontemporal
- |
  nontenured
- |
  nontheistic
- |
  nonthinking
- |
  nontoxic
- |
  nontrivial
- |
  nontropical
- |
  nontypical
- |
  nonunified
- |
  nonuniform
- |
  nonunion
- |
  nonuniversal
- |
  nonurban
- |
  nonuser
- |
  nonvascular
- |
  nonvenomous
- |
  nonverbal
- |
  nonviable
- |
  nonviolence
- |
  nonviolent
- |
  nonviolently
- |
  nonvirulent
- |
  nonvisual
- |
  nonvocal
- |
  nonvolatile
- |
  nonvolcanic
- |
  nonvoter
- |
  nonvoting
- |
  nonwhite
- |
  nonworker
- |
  nonworking
- |
  nonwoven
- |
  nonyielding
- |
  nonzero
- |
  noodle
- |
  noonday
- |
  noontide
- |
  noontime
- |
  noose
- |
  Nootka
- |
  noplace
- |
  Nordic
- |
  Noreen
- |
  Norfolk
- |
  Norgay
- |
  Norma
- |
  normal
- |
  normalcy
- |
  normalise
- |
  normality
- |
  normalize
- |
  normalizer
- |
  normally
- |
  Norman
- |
  Normandy
- |
  normative
- |
  normatively
- |
  Norplant
- |
  Norris
- |
  Norse
- |
  Norseman
- |
  North
- |
  north
- |
  Northampton
- |
  northbound
- |
  Northeast
- |
  northeast
- |
  northeaster
- |
  northeastern
- |
  norther
- |
  northerly
- |
  northern
- |
  Northerner
- |
  northerner
- |
  northernmost
- |
  Northumbria
- |
  Northumbrian
- |
  northward
- |
  northwardly
- |
  northwards
- |
  Northwest
- |
  northwest
- |
  northwestern
- |
  Norton
- |
  Norway
- |
  Norwegian
- |
  Norwich
- |
  nosebleed
- |
  nosecone
- |
  nosed
- |
  nosedive
- |
  nosedove
- |
  nosegay
- |
  nosepiece
- |
  nosey
- |
  nosher
- |
  nosily
- |
  nosiness
- |
  nosological
- |
  nosologist
- |
  nosology
- |
  nostalgia
- |
  nostalgic
- |
  nostalgist
- |
  Nostradamus
- |
  nostril
- |
  nostrum
- |
  notability
- |
  notable
- |
  notably
- |
  notarial
- |
  notarization
- |
  notarize
- |
  notary
- |
  notation
- |
  notch
- |
  notchback
- |
  notebook
- |
  noted
- |
  notepaper
- |
  notes
- |
  noteworthy
- |
  nothing
- |
  nothingness
- |
  notice
- |
  noticeable
- |
  noticeably
- |
  notification
- |
  notifier
- |
  notify
- |
  notion
- |
  notional
- |
  notionally
- |
  notions
- |
  notoriety
- |
  notorious
- |
  notoriously
- |
  Nottingham
- |
  Nouakchott
- |
  nougat
- |
  nought
- |
  Noumea
- |
  noumena
- |
  noumenal
- |
  noumenon
- |
  nourish
- |
  nourishing
- |
  nourishment
- |
  novae
- |
  novel
- |
  novelette
- |
  novelist
- |
  novelistic
- |
  novelization
- |
  novelize
- |
  novella
- |
  novelle
- |
  novelly
- |
  novelty
- |
  November
- |
  novena
- |
  Novgorod
- |
  novice
- |
  noviciate
- |
  novitiate
- |
  Novocain
- |
  Novocaine
- |
  Novokuznetsk
- |
  Novosibirsk
- |
  nowadays
- |
  noway
- |
  noways
- |
  nowhere
- |
  nowise
- |
  noxious
- |
  noxiously
- |
  noxiousness
- |
  noyade
- |
  Noyes
- |
  nozzle
- |
  nuance
- |
  nuanced
- |
  nubbin
- |
  nubbly
- |
  nubby
- |
  Nubia
- |
  Nubian
- |
  nubile
- |
  nubility
- |
  nuclear
- |
  nucleate
- |
  nucleation
- |
  nuclei
- |
  nucleic
- |
  nucleolar
- |
  nucleoli
- |
  nucleolus
- |
  nucleon
- |
  nucleonic
- |
  nucleonics
- |
  nucleotide
- |
  nucleus
- |
  nuclide
- |
  nuclidic
- |
  nudge
- |
  nudism
- |
  nudist
- |
  nudity
- |
  nudnick
- |
  nudnik
- |
  nugatory
- |
  nugget
- |
  nuisance
- |
  Nukualofa
- |
  nullifidian
- |
  nullifier
- |
  nullify
- |
  nullity
- |
  numbed
- |
  number
- |
  numberless
- |
  Numbers
- |
  numbers
- |
  numbly
- |
  numbness
- |
  numbskull
- |
  numen
- |
  numerable
- |
  numeracy
- |
  numeral
- |
  numerate
- |
  numeration
- |
  numerator
- |
  numeric
- |
  numerical
- |
  numerically
- |
  numerologist
- |
  numerology
- |
  numerous
- |
  numerously
- |
  numerousness
- |
  Numidia
- |
  Numidian
- |
  numina
- |
  numinous
- |
  numismatic
- |
  numismatics
- |
  numismatist
- |
  numskull
- |
  Nunavut
- |
  nuncio
- |
  nuncupative
- |
  nunnery
- |
  nuptial
- |
  nuptials
- |
  Nuremberg
- |
  Nureyev
- |
  Nurnberg
- |
  nurse
- |
  nursemaid
- |
  nurser
- |
  nursery
- |
  nurseryman
- |
  nursing
- |
  nursling
- |
  nurture
- |
  nurturer
- |
  nurturing
- |
  nutation
- |
  nutcracker
- |
  nuthatch
- |
  nutmeat
- |
  nutmeg
- |
  nutpick
- |
  nutria
- |
  nutrient
- |
  nutriment
- |
  nutrimental
- |
  nutrition
- |
  nutritional
- |
  nutritionist
- |
  nutritious
- |
  nutritiously
- |
  nutritive
- |
  nutshell
- |
  nuttily
- |
  nuttiness
- |
  nutty
- |
  nuzzle
- |
  nuzzler
- |
  Nyasa
- |
  Nyasaland
- |
  nyctalopia
- |
  nylon
- |
  nylons
- |
  nymph
- |
  nymphaea
- |
  nymphaeum
- |
  nymphal
- |
  nymphean
- |
  nymphet
- |
  nymphlike
- |
  nymphomania
- |
  nymphomaniac
- |
  nystagmic
- |
  nystagmus
- |
  oafish
- |
  oafishly
- |
  oafishness
- |
  oaken
- |
  Oakland
- |
  Oakley
- |
  oakum
- |
  oared
- |
  oarlock
- |
  oarsman
- |
  oarsmanship
- |
  oarswoman
- |
  oases
- |
  oasis
- |
  oatcake
- |
  oaten
- |
  Oates
- |
  oatmeal
- |
  Oaxaca
- |
  Obadiah
- |
  obbligati
- |
  obbligato
- |
  obduracy
- |
  obdurate
- |
  obdurately
- |
  obdurateness
- |
  obedience
- |
  obedient
- |
  obediently
- |
  obeisance
- |
  obeisant
- |
  obeli
- |
  obelisk
- |
  obelus
- |
  obese
- |
  obesely
- |
  obeseness
- |
  obesity
- |
  obeyer
- |
  obfuscate
- |
  obfuscation
- |
  obfuscatory
- |
  obituary
- |
  object
- |
  objectify
- |
  objection
- |
  objective
- |
  objectively
- |
  objectivism
- |
  objectivist
- |
  objectivity
- |
  objectivize
- |
  objector
- |
  objet
- |
  objurgate
- |
  objurgation
- |
  objurgator
- |
  objurgatory
- |
  oblate
- |
  oblately
- |
  oblateness
- |
  oblation
- |
  oblational
- |
  oblatory
- |
  obligate
- |
  obligati
- |
  obligation
- |
  obligato
- |
  obligator
- |
  obligatorily
- |
  obligatory
- |
  oblige
- |
  obliger
- |
  obliging
- |
  obligingly
- |
  obligingness
- |
  oblique
- |
  obliquely
- |
  obliqueness
- |
  obliquity
- |
  obliterate
- |
  obliteration
- |
  obliterative
- |
  obliterator
- |
  oblivion
- |
  oblivious
- |
  obliviously
- |
  oblong
- |
  obloquial
- |
  obloquious
- |
  obloquy
- |
  obnoxious
- |
  obnoxiously
- |
  oboist
- |
  obscene
- |
  obscenely
- |
  obscenity
- |
  obscurantism
- |
  obscurantist
- |
  obscure
- |
  obscurely
- |
  obscureness
- |
  obscurity
- |
  obsequies
- |
  obsequious
- |
  obsequiously
- |
  obsequy
- |
  observable
- |
  observably
- |
  observance
- |
  observant
- |
  observantly
- |
  observation
- |
  observatory
- |
  observe
- |
  observer
- |
  obsess
- |
  obsessed
- |
  obsession
- |
  obsessional
- |
  obsessive
- |
  obsessively
- |
  obsidian
- |
  obsolesce
- |
  obsolescence
- |
  obsolescent
- |
  obsolete
- |
  obsoletely
- |
  obsoleteness
- |
  obsoletism
- |
  obstacle
- |
  obstetric
- |
  obstetrical
- |
  obstetrician
- |
  obstetrics
- |
  obstinacy
- |
  obstinate
- |
  obstinately
- |
  obstreperous
- |
  obstruct
- |
  obstructer
- |
  obstruction
- |
  obstructive
- |
  obstructor
- |
  obtain
- |
  obtainable
- |
  obtainer
- |
  obtainment
- |
  obtrude
- |
  obtruder
- |
  obtrusion
- |
  obtrusive
- |
  obtrusively
- |
  obtuse
- |
  obtusely
- |
  obtuseness
- |
  obtusity
- |
  obverse
- |
  obversely
- |
  obviate
- |
  obviation
- |
  obviator
- |
  obvious
- |
  obviously
- |
  obviousness
- |
  ocarina
- |
  occasion
- |
  occasional
- |
  occasionally
- |
  Occident
- |
  occident
- |
  Occidental
- |
  occidental
- |
  occipita
- |
  occipital
- |
  occiput
- |
  occlude
- |
  occlusion
- |
  occlusive
- |
  occult
- |
  occultation
- |
  occultism
- |
  occultist
- |
  occultly
- |
  occultness
- |
  occupancy
- |
  occupant
- |
  occupation
- |
  occupational
- |
  occupied
- |
  occupier
- |
  occupy
- |
  occur
- |
  occurrence
- |
  Ocean
- |
  ocean
- |
  oceanaria
- |
  oceanarium
- |
  oceanfront
- |
  oceangoing
- |
  Oceania
- |
  Oceanian
- |
  oceanic
- |
  oceanography
- |
  oceanology
- |
  Oceanside
- |
  Oceanus
- |
  ocelot
- |
  ocher
- |
  ocherous
- |
  ochery
- |
  ochlocracy
- |
  ochlocrat
- |
  ochlocratic
- |
  ochre
- |
  ochreous
- |
  Ockham
- |
  octagon
- |
  octagonal
- |
  octahedra
- |
  octahedral
- |
  octahedron
- |
  octal
- |
  octane
- |
  Octans
- |
  octant
- |
  octantal
- |
  octave
- |
  Octavia
- |
  Octavian
- |
  Octavius
- |
  octavo
- |
  octet
- |
  octette
- |
  octillion
- |
  octillionth
- |
  October
- |
  octogenarian
- |
  octopi
- |
  octopus
- |
  octosyllabic
- |
  octuplet
- |
  ocular
- |
  oculist
- |
  odalisk
- |
  odalisque
- |
  oddball
- |
  oddity
- |
  oddly
- |
  oddment
- |
  oddness
- |
  Odense
- |
  odeon
- |
  Odessa
- |
  Odets
- |
  odeum
- |
  odious
- |
  odiously
- |
  odiousness
- |
  odium
- |
  odometer
- |
  odontologist
- |
  odontology
- |
  odored
- |
  odoriferous
- |
  odorless
- |
  odorlessly
- |
  odorous
- |
  odorously
- |
  odorousness
- |
  odour
- |
  Odyssean
- |
  Odysseus
- |
  Odyssey
- |
  odyssey
- |
  oecumenical
- |
  oedema
- |
  Oedipal
- |
  oedipal
- |
  Oedipus
- |
  oenologist
- |
  oenology
- |
  oenophile
- |
  oenophilist
- |
  oesophagus
- |
  oestrogen
- |
  oestrous
- |
  oestrus
- |
  oeuvre
- |
  offal
- |
  offbeat
- |
  Offenbach
- |
  offence
- |
  offend
- |
  offended
- |
  offender
- |
  offending
- |
  offense
- |
  offensive
- |
  offensively
- |
  offer
- |
  offerer
- |
  offering
- |
  offeror
- |
  Offertory
- |
  offertory
- |
  offhand
- |
  offhanded
- |
  offhandedly
- |
  office
- |
  officeholder
- |
  officer
- |
  offices
- |
  official
- |
  officialdom
- |
  officialism
- |
  officially
- |
  officiant
- |
  officiate
- |
  officiation
- |
  officiator
- |
  officious
- |
  officiously
- |
  offing
- |
  offish
- |
  offishly
- |
  offishness
- |
  offkey
- |
  offline
- |
  offload
- |
  offprint
- |
  offscreen
- |
  offset
- |
  offshoot
- |
  offshore
- |
  offside
- |
  offsides
- |
  offspring
- |
  offstage
- |
  offtrack
- |
  often
- |
  oftentimes
- |
  ofttimes
- |
  Ogbomosho
- |
  ogeed
- |
  ogival
- |
  ogive
- |
  Oglala
- |
  ogler
- |
  Oglethorpe
- |
  ogreish
- |
  ogress
- |
  ogrish
- |
  Ohioan
- |
  ohmic
- |
  ohmmeter
- |
  oilcloth
- |
  oiled
- |
  oiler
- |
  oilfield
- |
  oilily
- |
  oiliness
- |
  oilskin
- |
  oilskins
- |
  ointment
- |
  Ojibwa
- |
  Ojibway
- |
  Okavango
- |
  Okayama
- |
  Okeechobee
- |
  Okefenokee
- |
  Okhotsk
- |
  Okinawa
- |
  Okinawan
- |
  Oklahoma
- |
  Oklahoman
- |
  olden
- |
  Oldham
- |
  oldie
- |
  oldish
- |
  oldness
- |
  oldster
- |
  Olduvai
- |
  oleaginous
- |
  oleander
- |
  oleomargarin
- |
  olestra
- |
  olfaction
- |
  olfactory
- |
  oligarch
- |
  oligarchic
- |
  oligarchical
- |
  oligarchy
- |
  Oligocene
- |
  oligopolist
- |
  oligopoly
- |
  Olive
- |
  olive
- |
  Oliver
- |
  Olives
- |
  Olivet
- |
  Olivia
- |
  Olivier
- |
  olivine
- |
  Ollie
- |
  Olmec
- |
  Olmsted
- |
  Olympia
- |
  Olympiad
- |
  Olympian
- |
  Olympic
- |
  Olympics
- |
  Olympus
- |
  Omagh
- |
  Omaha
- |
  Omani
- |
  ombudsman
- |
  Omdurman
- |
  omega
- |
  omelet
- |
  omelette
- |
  omicron
- |
  omikron
- |
  ominous
- |
  ominously
- |
  ominousness
- |
  omissible
- |
  omission
- |
  omnibus
- |
  omnipotence
- |
  Omnipotent
- |
  omnipotent
- |
  omnipotently
- |
  omnipresence
- |
  omnipresent
- |
  omniscience
- |
  Omniscient
- |
  omniscient
- |
  omnisciently
- |
  omnivore
- |
  omnivorous
- |
  omnivorously
- |
  omphaloi
- |
  omphalos
- |
  onanism
- |
  onanist
- |
  onanistic
- |
  Onassis
- |
  oncogene
- |
  oncogenesis
- |
  oncogenic
- |
  oncogenicity
- |
  oncologic
- |
  oncological
- |
  oncologist
- |
  oncology
- |
  oncoming
- |
  Oneida
- |
  oneiric
- |
  oneiromancy
- |
  oneness
- |
  onerous
- |
  onerously
- |
  onerousness
- |
  oneself
- |
  onetime
- |
  ongoing
- |
  onion
- |
  onionskin
- |
  online
- |
  onlooker
- |
  onlooking
- |
  onomasiology
- |
  onomatopoeia
- |
  onomatopoeic
- |
  Onondaga
- |
  Onondagan
- |
  onrush
- |
  onrushing
- |
  onscreen
- |
  onset
- |
  onshore
- |
  onslaught
- |
  onstage
- |
  Ontarian
- |
  Ontario
- |
  ontic
- |
  ontogenetic
- |
  ontogenic
- |
  ontogeny
- |
  ontological
- |
  ontologist
- |
  ontology
- |
  onward
- |
  onwards
- |
  oocyte
- |
  oodles
- |
  oogenesis
- |
  oogenetic
- |
  oogonia
- |
  oogonium
- |
  oolite
- |
  oolitic
- |
  oologic
- |
  oological
- |
  oologically
- |
  oologist
- |
  oology
- |
  oomph
- |
  ooziness
- |
  opacity
- |
  opalesce
- |
  opalescence
- |
  opalescent
- |
  opaline
- |
  opaque
- |
  opaquely
- |
  opaqueness
- |
  opener
- |
  openhanded
- |
  openhandedly
- |
  opening
- |
  openly
- |
  openness
- |
  openwork
- |
  opera
- |
  operability
- |
  operable
- |
  operably
- |
  operand
- |
  operant
- |
  operate
- |
  operatic
- |
  operatically
- |
  operating
- |
  operation
- |
  operational
- |
  operative
- |
  operatively
- |
  operator
- |
  operetta
- |
  operose
- |
  Ophelia
- |
  Ophiuchus
- |
  ophthalmic
- |
  opiate
- |
  opine
- |
  opinion
- |
  opinionated
- |
  opium
- |
  Oporto
- |
  opossum
- |
  Oppenheimer
- |
  opponent
- |
  opportune
- |
  opportunely
- |
  opportunism
- |
  opportunist
- |
  opportunity
- |
  opposability
- |
  opposable
- |
  oppose
- |
  opposed
- |
  opposer
- |
  opposing
- |
  opposite
- |
  oppositely
- |
  oppositeness
- |
  opposition
- |
  oppositional
- |
  oppress
- |
  oppressed
- |
  oppression
- |
  oppressive
- |
  oppressively
- |
  oppressor
- |
  opprobrious
- |
  opprobrium
- |
  optic
- |
  optical
- |
  optically
- |
  optician
- |
  optics
- |
  optima
- |
  optimal
- |
  optimality
- |
  optimally
- |
  optimism
- |
  optimist
- |
  optimistic
- |
  optimization
- |
  optimize
- |
  optimum
- |
  option
- |
  optional
- |
  optionality
- |
  optionally
- |
  optometric
- |
  optometrist
- |
  optometry
- |
  opulence
- |
  opulent
- |
  opulently
- |
  oracle
- |
  oracular
- |
  oracularity
- |
  oracularly
- |
  orally
- |
  orang
- |
  Orange
- |
  orange
- |
  orangeade
- |
  orangery
- |
  orangutan
- |
  orangutang
- |
  Oranjestad
- |
  orate
- |
  oration
- |
  orator
- |
  oratorical
- |
  oratorically
- |
  oratorio
- |
  oratory
- |
  orbicular
- |
  orbicularity
- |
  orbicularly
- |
  orbit
- |
  orbital
- |
  orbiter
- |
  orchard
- |
  orchardist
- |
  orchestra
- |
  orchestral
- |
  orchestrally
- |
  orchestrate
- |
  orchestrator
- |
  orchid
- |
  ordain
- |
  ordainer
- |
  ordainment
- |
  ordeal
- |
  order
- |
  orderer
- |
  orderliness
- |
  orderly
- |
  orders
- |
  ordinal
- |
  ordinance
- |
  ordinarily
- |
  ordinariness
- |
  ordinary
- |
  ordinate
- |
  ordination
- |
  ordines
- |
  ordnance
- |
  ordonnance
- |
  Ordovician
- |
  ordure
- |
  oread
- |
  oregano
- |
  Oregon
- |
  Oregonian
- |
  Orenburg
- |
  Orestes
- |
  organ
- |
  organdie
- |
  organdy
- |
  organelle
- |
  organic
- |
  organically
- |
  organicity
- |
  organisation
- |
  organise
- |
  organised
- |
  organiser
- |
  organism
- |
  organismic
- |
  organist
- |
  organization
- |
  organize
- |
  organized
- |
  organizer
- |
  organon
- |
  organza
- |
  orgasm
- |
  orgasmic
- |
  orgasmically
- |
  orgastic
- |
  orgastically
- |
  orgiast
- |
  orgiastic
- |
  orgulous
- |
  oriel
- |
  Orient
- |
  orient
- |
  Oriental
- |
  oriental
- |
  Orientalism
- |
  Orientalist
- |
  orientalize
- |
  orientally
- |
  orientate
- |
  orientation
- |
  oriented
- |
  orienteer
- |
  orienteering
- |
  orifice
- |
  orificial
- |
  oriflamme
- |
  origami
- |
  origin
- |
  original
- |
  originality
- |
  originally
- |
  originate
- |
  origination
- |
  originator
- |
  origins
- |
  Orinoco
- |
  oriole
- |
  Orion
- |
  orison
- |
  Orkney
- |
  Orlando
- |
  Orleans
- |
  Orlon
- |
  Ormazd
- |
  ormolu
- |
  Ormuz
- |
  ornament
- |
  ornamental
- |
  ornamentally
- |
  ornate
- |
  ornately
- |
  ornateness
- |
  orneriness
- |
  ornery
- |
  ornithologic
- |
  ornithology
- |
  orogenesis
- |
  orogenic
- |
  orogeny
- |
  orographic
- |
  orographical
- |
  orography
- |
  orotund
- |
  orotundity
- |
  orphan
- |
  orphanage
- |
  orphanhood
- |
  Orpheus
- |
  Orphic
- |
  Orphism
- |
  orrery
- |
  Orrin
- |
  orris
- |
  Orson
- |
  orthodontia
- |
  orthodontic
- |
  orthodontics
- |
  orthodontist
- |
  orthodonture
- |
  Orthodox
- |
  orthodox
- |
  orthodoxly
- |
  orthodoxy
- |
  orthogonal
- |
  orthogonally
- |
  orthographic
- |
  orthography
- |
  orthopaedic
- |
  orthopaedics
- |
  orthopaedist
- |
  orthopedic
- |
  orthopedics
- |
  orthopedist
- |
  orthoses
- |
  orthosis
- |
  orthotic
- |
  orthotics
- |
  orthotist
- |
  Orval
- |
  Orville
- |
  Orwell
- |
  Orwellian
- |
  Osage
- |
  Osaka
- |
  Oscar
- |
  Osceola
- |
  oscillate
- |
  oscillation
- |
  oscillator
- |
  oscillatory
- |
  oscilloscope
- |
  oscitancy
- |
  oscitation
- |
  osculant
- |
  osculate
- |
  osculation
- |
  osculatory
- |
  Oshawa
- |
  Oshkosh
- |
  osier
- |
  Osiris
- |
  Osman
- |
  osmic
- |
  osmically
- |
  osmium
- |
  osmose
- |
  osmosis
- |
  osmotic
- |
  osmotically
- |
  osprey
- |
  osseous
- |
  ossific
- |
  ossification
- |
  ossify
- |
  ossuary
- |
  osteitis
- |
  ostensible
- |
  ostensibly
- |
  ostensive
- |
  ostentation
- |
  ostentatious
- |
  osteopath
- |
  osteopathic
- |
  osteopathy
- |
  osteoporoses
- |
  osteoporosis
- |
  osteoporotic
- |
  Ostia
- |
  ostler
- |
  ostmark
- |
  ostomy
- |
  ostracism
- |
  ostracize
- |
  Ostrava
- |
  ostrich
- |
  Ostrogoth
- |
  Oswald
- |
  Othello
- |
  other
- |
  others
- |
  otherwise
- |
  otherworld
- |
  otherworldly
- |
  Othman
- |
  otiose
- |
  otiosely
- |
  otitis
- |
  Ottawa
- |
  otter
- |
  Ottoman
- |
  ottoman
- |
  Ouagadougou
- |
  oubliette
- |
  ought
- |
  ouguiya
- |
  Ouija
- |
  Oujda
- |
  ounce
- |
  ourself
- |
  ourselves
- |
  ouster
- |
  ousting
- |
  outage
- |
  outargue
- |
  outback
- |
  outbalance
- |
  outbargain
- |
  outbid
- |
  outboard
- |
  outboast
- |
  outbound
- |
  outbreak
- |
  outbuilding
- |
  outburst
- |
  outcast
- |
  outclass
- |
  outcome
- |
  outcrop
- |
  outcropping
- |
  outcry
- |
  outdated
- |
  outdid
- |
  outdistance
- |
  outdo
- |
  outdone
- |
  outdoor
- |
  outdoors
- |
  outdraw
- |
  outdrawn
- |
  outdrew
- |
  outearn
- |
  outer
- |
  outermost
- |
  outerwear
- |
  outface
- |
  outfall
- |
  outfield
- |
  outfielder
- |
  outfight
- |
  outfit
- |
  outfitter
- |
  outflank
- |
  outflatter
- |
  outflow
- |
  outfought
- |
  outfox
- |
  outgo
- |
  outgoing
- |
  outgrew
- |
  outgrow
- |
  outgrown
- |
  outgrowth
- |
  outguess
- |
  outgun
- |
  outhit
- |
  outhouse
- |
  outing
- |
  outland
- |
  outlander
- |
  outlandish
- |
  outlandishly
- |
  outlands
- |
  outlast
- |
  outlaw
- |
  outlawry
- |
  outlay
- |
  outlet
- |
  outline
- |
  outlive
- |
  outlook
- |
  outlying
- |
  outmaneuver
- |
  outmanoeuvre
- |
  outmatch
- |
  outmoded
- |
  outnumber
- |
  outpace
- |
  outpatient
- |
  outperform
- |
  outplacement
- |
  outplay
- |
  outpoint
- |
  outpost
- |
  outpouring
- |
  outproduce
- |
  outpull
- |
  output
- |
  outrace
- |
  outrage
- |
  outraged
- |
  outrageous
- |
  outrageously
- |
  outran
- |
  outrank
- |
  outre
- |
  outreach
- |
  outreason
- |
  outrider
- |
  outrigger
- |
  outright
- |
  outrun
- |
  outscore
- |
  outsell
- |
  outset
- |
  outshine
- |
  outshone
- |
  outshout
- |
  outside
- |
  outsider
- |
  outsize
- |
  outsized
- |
  outskirt
- |
  outskirts
- |
  outsmart
- |
  outsold
- |
  outsource
- |
  outsourcing
- |
  outspend
- |
  outspoken
- |
  outspokenly
- |
  outspread
- |
  outstanding
- |
  outstation
- |
  outstay
- |
  outstretch
- |
  outstretched
- |
  outstrip
- |
  outtake
- |
  outvote
- |
  outwait
- |
  outwalk
- |
  outward
- |
  outwardly
- |
  outwards
- |
  outwear
- |
  outweigh
- |
  outwit
- |
  outwore
- |
  outwork
- |
  outworn
- |
  outyell
- |
  ovarian
- |
  ovary
- |
  ovate
- |
  ovately
- |
  ovation
- |
  ovenbird
- |
  overabundant
- |
  overachieve
- |
  overachiever
- |
  overact
- |
  overactive
- |
  overage
- |
  overall
- |
  overalls
- |
  overambition
- |
  overanalyze
- |
  overanxious
- |
  overarching
- |
  overarm
- |
  overassured
- |
  overate
- |
  overattached
- |
  overawe
- |
  overawed
- |
  overbalance
- |
  overbear
- |
  overbearing
- |
  overbid
- |
  overbite
- |
  overblown
- |
  overboard
- |
  overbold
- |
  overbook
- |
  overbought
- |
  overbuild
- |
  overburden
- |
  overburdened
- |
  overbuy
- |
  overcame
- |
  overcapacity
- |
  overcareful
- |
  overcast
- |
  overcautious
- |
  overcharge
- |
  overcharging
- |
  overclothes
- |
  overcloud
- |
  overcoat
- |
  overcome
- |
  overconcern
- |
  overcook
- |
  overcool
- |
  overcritical
- |
  overcrowd
- |
  overcrowded
- |
  overcrowding
- |
  overcurious
- |
  overdecorate
- |
  overdesirous
- |
  overdetailed
- |
  overdevelop
- |
  overdid
- |
  overdo
- |
  overdone
- |
  overdose
- |
  overdraft
- |
  overdraw
- |
  overdrawn
- |
  overdress
- |
  overdrew
- |
  overdrive
- |
  overdub
- |
  overdue
- |
  overeager
- |
  overeat
- |
  overeaten
- |
  overeater
- |
  overeating
- |
  overeducate
- |
  overeducated
- |
  overemphasis
- |
  overemphatic
- |
  overendowed
- |
  overestimate
- |
  overexcite
- |
  overexcited
- |
  overexercise
- |
  overexert
- |
  overexertion
- |
  overexpand
- |
  overexplicit
- |
  overexpose
- |
  overexposure
- |
  overextend
- |
  overextended
- |
  overfamiliar
- |
  overfanciful
- |
  overfatigued
- |
  overfed
- |
  overfeed
- |
  overfill
- |
  overflew
- |
  overflight
- |
  overflow
- |
  overflown
- |
  overfly
- |
  overfond
- |
  overfull
- |
  overgenerous
- |
  overgraze
- |
  overgrew
- |
  overgrow
- |
  overgrown
- |
  overgrowth
- |
  overhand
- |
  overhanded
- |
  overhang
- |
  overhastily
- |
  overhasty
- |
  overhaul
- |
  overhead
- |
  overheads
- |
  overhear
- |
  overheard
- |
  overheat
- |
  overheated
- |
  overhung
- |
  overhurried
- |
  overimpress
- |
  overincline
- |
  overindulge
- |
  overinflate
- |
  overinsure
- |
  overintense
- |
  overinterest
- |
  overinvest
- |
  overjoy
- |
  overjoyed
- |
  overkill
- |
  overlaid
- |
  overlain
- |
  overland
- |
  overlap
- |
  overlarge
- |
  overlavish
- |
  overlay
- |
  overleaf
- |
  overleap
- |
  overleapt
- |
  overlearn
- |
  overlie
- |
  overload
- |
  overloaded
- |
  overlong
- |
  overlook
- |
  overlord
- |
  overly
- |
  overmagnify
- |
  overmaster
- |
  overmatch
- |
  overmedicate
- |
  overmodest
- |
  overmodify
- |
  overmuch
- |
  overnice
- |
  overnight
- |
  overoptimism
- |
  overpaid
- |
  overpass
- |
  overpay
- |
  overplay
- |
  overpopulate
- |
  overpower
- |
  overpowerful
- |
  overpowering
- |
  overpraise
- |
  overprecise
- |
  overprice
- |
  overpriced
- |
  overprint
- |
  overproduce
- |
  overprompt
- |
  overprotect
- |
  overproud
- |
  overran
- |
  overrate
- |
  overrated
- |
  overreach
- |
  overreacher
- |
  overreaching
- |
  overreact
- |
  overreaction
- |
  overrefine
- |
  overrefined
- |
  overregulate
- |
  overridden
- |
  override
- |
  overriding
- |
  overridingly
- |
  overrigid
- |
  overripe
- |
  overripen
- |
  overroast
- |
  overrode
- |
  overrule
- |
  overrun
- |
  oversalt
- |
  oversaw
- |
  overscale
- |
  overscaled
- |
  oversea
- |
  overseas
- |
  oversee
- |
  overseen
- |
  overseer
- |
  oversell
- |
  oversevere
- |
  oversexed
- |
  overshadow
- |
  oversharp
- |
  overshoe
- |
  overshoot
- |
  overshot
- |
  oversight
- |
  oversimple
- |
  oversimplify
- |
  oversize
- |
  oversized
- |
  overskirt
- |
  oversleep
- |
  overslept
- |
  oversold
- |
  overspend
- |
  overspent
- |
  overspill
- |
  overspread
- |
  overstaff
- |
  overstate
- |
  overstay
- |
  oversteer
- |
  overstep
- |
  overstock
- |
  overstrain
- |
  overstress
- |
  overstretch
- |
  overstrict
- |
  overstrung
- |
  overstuff
- |
  overstuffed
- |
  oversubtle
- |
  oversupply
- |
  overt
- |
  overtake
- |
  overtaken
- |
  overtax
- |
  overtaxation
- |
  overthrew
- |
  overthrow
- |
  overthrown
- |
  overtime
- |
  overtire
- |
  overtired
- |
  overtly
- |
  overtness
- |
  overtone
- |
  overtones
- |
  overtook
- |
  overtop
- |
  overtrain
- |
  overtrick
- |
  overture
- |
  overtures
- |
  overturn
- |
  overuse
- |
  overvalue
- |
  overvalued
- |
  overview
- |
  overviolent
- |
  overweary
- |
  overweening
- |
  overweigh
- |
  overweight
- |
  overwhelm
- |
  overwhelmed
- |
  overwhelming
- |
  overwilling
- |
  overwind
- |
  overwinter
- |
  overwork
- |
  overworked
- |
  overwritten
- |
  overwrought
- |
  overzealous
- |
  oviduct
- |
  Oviedo
- |
  ovine
- |
  oviparity
- |
  oviparous
- |
  ovoid
- |
  ovoidal
- |
  ovular
- |
  ovulate
- |
  ovulation
- |
  ovulatory
- |
  ovule
- |
  Owens
- |
  owing
- |
  owlet
- |
  owlish
- |
  owlishly
- |
  owned
- |
  owner
- |
  ownership
- |
  oxblood
- |
  oxbow
- |
  Oxbridge
- |
  Oxford
- |
  oxford
- |
  Oxfordshire
- |
  oxidant
- |
  oxidation
- |
  oxidative
- |
  oxidatively
- |
  oxide
- |
  oxidic
- |
  oxidise
- |
  oxidizable
- |
  oxidization
- |
  oxidize
- |
  oxidizer
- |
  Oxnard
- |
  Oxonian
- |
  oxyacetylene
- |
  oxygen
- |
  oxygenate
- |
  oxygenation
- |
  oxygenic
- |
  oxygenous
- |
  oxymora
- |
  oxymoron
- |
  oxymoronic
- |
  oyster
- |
  oystering
- |
  oysterman
- |
  Ozarks
- |
  ozone
- |
  ozonic
- |
  ozonosphere
- |
  Pablum
- |
  pabulum
- |
  pacemaker
- |
  pacemaking
- |
  pacer
- |
  pacesetter
- |
  Pachuca
- |
  pachyderm
- |
  pachydermal
- |
  pachydermous
- |
  pachysandra
- |
  Pacific
- |
  pacific
- |
  pacifically
- |
  pacification
- |
  pacificatory
- |
  pacifier
- |
  pacifism
- |
  pacifist
- |
  pacifistic
- |
  pacify
- |
  package
- |
  packager
- |
  packaging
- |
  packed
- |
  packer
- |
  packet
- |
  packetboat
- |
  packhorse
- |
  packing
- |
  packinghouse
- |
  packsaddle
- |
  packthread
- |
  Padang
- |
  padded
- |
  padding
- |
  paddle
- |
  paddleboard
- |
  paddler
- |
  paddock
- |
  paddy
- |
  Paderewski
- |
  padlock
- |
  Padre
- |
  padre
- |
  padrone
- |
  Padua
- |
  paean
- |
  paediatric
- |
  paediatrics
- |
  paedophile
- |
  paella
- |
  Paestum
- |
  pagan
- |
  Paganini
- |
  paganish
- |
  paganism
- |
  paganize
- |
  pageant
- |
  pageantry
- |
  pageboy
- |
  pager
- |
  paginate
- |
  pagination
- |
  pagoda
- |
  Pahlavi
- |
  pailful
- |
  Paine
- |
  pained
- |
  painful
- |
  painfully
- |
  painkiller
- |
  painkilling
- |
  painless
- |
  painlessly
- |
  painlessness
- |
  pains
- |
  painstaking
- |
  paint
- |
  paintbox
- |
  paintbrush
- |
  painter
- |
  painting
- |
  paints
- |
  pairing
- |
  paisa
- |
  paisley
- |
  Paiute
- |
  pajamas
- |
  Pakistan
- |
  Pakistani
- |
  palace
- |
  paladin
- |
  palaestra
- |
  palaestrae
- |
  palanquin
- |
  palatability
- |
  palatable
- |
  palatably
- |
  palatal
- |
  palatalize
- |
  palate
- |
  palatial
- |
  palatially
- |
  palatinate
- |
  palatine
- |
  Palau
- |
  palaver
- |
  Palawan
- |
  paleface
- |
  palely
- |
  Palembang
- |
  paleness
- |
  paleobiology
- |
  Paleocene
- |
  paleographer
- |
  paleographic
- |
  paleography
- |
  Paleolithic
- |
  paleolithic
- |
  paleontology
- |
  Paleozoic
- |
  Palermo
- |
  Palestine
- |
  Palestinian
- |
  palette
- |
  palfrey
- |
  palimony
- |
  palimpsest
- |
  palimpsestic
- |
  palindrome
- |
  palindromic
- |
  palindromist
- |
  paling
- |
  palingenesis
- |
  palingenetic
- |
  palisade
- |
  palisaded
- |
  Palisades
- |
  palisades
- |
  palish
- |
  Palladian
- |
  Palladio
- |
  palladium
- |
  pallbearer
- |
  pallet
- |
  pallia
- |
  palliate
- |
  palliation
- |
  palliative
- |
  palliator
- |
  pallid
- |
  pallidly
- |
  pallidness
- |
  pallium
- |
  pallor
- |
  Palma
- |
  palmate
- |
  palmated
- |
  palmately
- |
  Palmer
- |
  Palmerston
- |
  palmetto
- |
  palmist
- |
  palmistry
- |
  palmtop
- |
  palmy
- |
  Palomar
- |
  palomino
- |
  palpability
- |
  palpable
- |
  palpably
- |
  palpate
- |
  palpation
- |
  palpitate
- |
  palpitating
- |
  palpitation
- |
  palpitations
- |
  palsied
- |
  palsy
- |
  palter
- |
  paltriness
- |
  paltry
- |
  paludal
- |
  Pamela
- |
  Pamir
- |
  Pamirs
- |
  Pamlico
- |
  Pampa
- |
  pampa
- |
  pampas
- |
  pamper
- |
  pamphlet
- |
  pamphleteer
- |
  Pamplona
- |
  panacea
- |
  panacean
- |
  panache
- |
  Panama
- |
  panama
- |
  Panamanian
- |
  panatela
- |
  Panay
- |
  pancake
- |
  Panchiao
- |
  panchromatic
- |
  pancreas
- |
  pancreatic
- |
  pancreatitis
- |
  panda
- |
  pandect
- |
  pandectist
- |
  pandemic
- |
  pandemonium
- |
  pander
- |
  panderer
- |
  Pandora
- |
  pandowdy
- |
  panegyric
- |
  panegyrical
- |
  panegyrist
- |
  panel
- |
  paneled
- |
  paneling
- |
  panelist
- |
  panelled
- |
  panelling
- |
  panful
- |
  Pangaea
- |
  panhandle
- |
  panhandler
- |
  panic
- |
  panicky
- |
  panicle
- |
  panicled
- |
  panier
- |
  Panjabi
- |
  panjandra
- |
  panjandrum
- |
  Pankhurst
- |
  pannier
- |
  panocha
- |
  panoplied
- |
  panoply
- |
  panorama
- |
  panoramic
- |
  panpipe
- |
  pansy
- |
  pantaloon
- |
  pantaloons
- |
  pantheism
- |
  pantheist
- |
  pantheistic
- |
  pantheon
- |
  panther
- |
  pantie
- |
  panties
- |
  pantingly
- |
  pantomime
- |
  pantomimic
- |
  pantomimist
- |
  pantry
- |
  pants
- |
  pantsuit
- |
  panty
- |
  pantyhose
- |
  pantyliner
- |
  pantywaist
- |
  Papacy
- |
  papacy
- |
  Papago
- |
  papain
- |
  papal
- |
  papally
- |
  Papandreou
- |
  paparazzi
- |
  paparazzo
- |
  papaw
- |
  papaya
- |
  Papeete
- |
  paper
- |
  paperback
- |
  paperboard
- |
  paperbound
- |
  paperboy
- |
  paperer
- |
  papergirl
- |
  paperhanger
- |
  paperhanging
- |
  paperless
- |
  papers
- |
  paperweight
- |
  paperwork
- |
  papery
- |
  papilla
- |
  papillae
- |
  papillary
- |
  papism
- |
  papist
- |
  papistical
- |
  papistry
- |
  papoose
- |
  paprika
- |
  Papuan
- |
  papular
- |
  papule
- |
  papyri
- |
  papyrus
- |
  parable
- |
  parabola
- |
  parabolae
- |
  parabolic
- |
  Paracelsus
- |
  parachronism
- |
  parachute
- |
  parachutist
- |
  parade
- |
  parader
- |
  paradigm
- |
  paradigmatic
- |
  paradisaic
- |
  paradisaical
- |
  Paradise
- |
  paradise
- |
  paradisiac
- |
  paradisiacal
- |
  paradox
- |
  paradoxical
- |
  paraffin
- |
  paraffine
- |
  paraffinic
- |
  parafoil
- |
  paraglider
- |
  paragon
- |
  paragraph
- |
  Paraguay
- |
  Paraguayan
- |
  Paraiba
- |
  parakeet
- |
  paralegal
- |
  parallactic
- |
  parallax
- |
  parallel
- |
  parallelism
- |
  parallepiped
- |
  paralogism
- |
  paralogist
- |
  paralyse
- |
  paralysed
- |
  paralyses
- |
  paralysing
- |
  paralysis
- |
  paralytic
- |
  paralyze
- |
  paralyzed
- |
  paralyzing
- |
  paralyzingly
- |
  Paramaribo
- |
  paramecia
- |
  paramecium
- |
  paramedic
- |
  paramedical
- |
  parameter
- |
  parameters
- |
  parametric
- |
  paramilitary
- |
  paramount
- |
  paramour
- |
  Parana
- |
  paranoia
- |
  paranoiac
- |
  paranoic
- |
  paranoically
- |
  paranoid
- |
  paranormal
- |
  paranormally
- |
  parapet
- |
  parapeted
- |
  paraphilia
- |
  paraphiliac
- |
  paraphrase
- |
  paraphraser
- |
  paraphrasis
- |
  paraphrastic
- |
  paraplegia
- |
  paraplegic
- |
  paraquat
- |
  parasite
- |
  parasitic
- |
  parasitical
- |
  parasitism
- |
  parasitize
- |
  parasitology
- |
  parasol
- |
  paratactic
- |
  parataxis
- |
  parathion
- |
  parathyroid
- |
  paratrooper
- |
  paratroops
- |
  paratyphoid
- |
  parboil
- |
  parcel
- |
  parch
- |
  parched
- |
  parchment
- |
  pardon
- |
  pardonable
- |
  pardonably
- |
  pardoner
- |
  paregoric
- |
  parent
- |
  parentage
- |
  parental
- |
  parentheses
- |
  parenthesis
- |
  parenthesize
- |
  parenthetic
- |
  parenthood
- |
  parenting
- |
  parer
- |
  pareses
- |
  paresis
- |
  paretic
- |
  pareve
- |
  parfait
- |
  parhelia
- |
  parhelion
- |
  pariah
- |
  Parian
- |
  Paricutin
- |
  parietal
- |
  parietals
- |
  parimutuel
- |
  paring
- |
  Paris
- |
  parish
- |
  parishioner
- |
  Parisian
- |
  parity
- |
  parka
- |
  parked
- |
  Parker
- |
  parking
- |
  Parkinson
- |
  Parkinsonism
- |
  parkland
- |
  Parkman
- |
  Parks
- |
  parkway
- |
  parlance
- |
  parlay
- |
  parley
- |
  Parliament
- |
  parliament
- |
  parlor
- |
  parlour
- |
  parlous
- |
  parlously
- |
  parlousness
- |
  Parma
- |
  Parmenides
- |
  Parmesan
- |
  parmigiana
- |
  parmigiano
- |
  Parnaiba
- |
  Parnassian
- |
  Parnassus
- |
  Parnell
- |
  parochial
- |
  parochialism
- |
  parochiality
- |
  parochially
- |
  parodic
- |
  parodist
- |
  parody
- |
  parole
- |
  parolee
- |
  paronomasia
- |
  paronym
- |
  paronymic
- |
  paronymous
- |
  paronymy
- |
  Paros
- |
  paroxysm
- |
  paroxysmal
- |
  parquet
- |
  parquetry
- |
  parrakeet
- |
  Parramatta
- |
  parricidal
- |
  parricide
- |
  Parrish
- |
  parrot
- |
  parry
- |
  parse
- |
  parsec
- |
  parser
- |
  parsimonious
- |
  parsimony
- |
  parsley
- |
  parsnip
- |
  parson
- |
  parsonage
- |
  partake
- |
  partaken
- |
  partaker
- |
  parted
- |
  parterre
- |
  Parthenon
- |
  Parthia
- |
  Parthian
- |
  partial
- |
  partiality
- |
  partially
- |
  partialness
- |
  participant
- |
  participate
- |
  participator
- |
  participial
- |
  participle
- |
  particle
- |
  particolored
- |
  particular
- |
  particularly
- |
  particulate
- |
  particulates
- |
  parting
- |
  partisan
- |
  partisanship
- |
  partite
- |
  partition
- |
  partitioned
- |
  partitive
- |
  partizan
- |
  partly
- |
  partner
- |
  partnership
- |
  partook
- |
  partridge
- |
  parts
- |
  parturient
- |
  parturition
- |
  partway
- |
  party
- |
  parve
- |
  parvenu
- |
  Pasadena
- |
  PASCAL
- |
  Pascal
- |
  pascal
- |
  paschal
- |
  pasha
- |
  Pashto
- |
  pasquinade
- |
  passable
- |
  passably
- |
  passage
- |
  passageway
- |
  passbook
- |
  passe
- |
  passel
- |
  passenger
- |
  passer
- |
  passerby
- |
  passerine
- |
  passersby
- |
  passim
- |
  passing
- |
  passingly
- |
  Passion
- |
  passion
- |
  passionate
- |
  passionately
- |
  passionless
- |
  passivate
- |
  passive
- |
  passively
- |
  passiveness
- |
  passivity
- |
  passkey
- |
  Passover
- |
  passport
- |
  password
- |
  pasta
- |
  paste
- |
  pasteboard
- |
  pastel
- |
  pastern
- |
  Pasternak
- |
  Pasteur
- |
  Pasteurian
- |
  pasteurize
- |
  pasteurizer
- |
  pastiche
- |
  pastil
- |
  pastille
- |
  pastime
- |
  pastiness
- |
  pastor
- |
  pastoral
- |
  pastorale
- |
  pastorali
- |
  pastoralism
- |
  pastoralist
- |
  pastorally
- |
  pastorate
- |
  pastrami
- |
  pastry
- |
  pasturage
- |
  pasture
- |
  pasty
- |
  pataca
- |
  Patagonia
- |
  Patagonian
- |
  patch
- |
  patchily
- |
  patchiness
- |
  patchwork
- |
  patchy
- |
  patella
- |
  patellae
- |
  patellar
- |
  paten
- |
  patent
- |
  patentable
- |
  patentee
- |
  patently
- |
  paternal
- |
  paternalism
- |
  paternalist
- |
  paternally
- |
  paternity
- |
  Paternoster
- |
  paternoster
- |
  Paterson
- |
  pathbreaking
- |
  pathetic
- |
  pathetically
- |
  pathfinder
- |
  pathless
- |
  pathname
- |
  pathogen
- |
  pathogenesis
- |
  pathogenic
- |
  pathogenous
- |
  pathologic
- |
  pathological
- |
  pathologist
- |
  pathology
- |
  pathos
- |
  pathway
- |
  patience
- |
  patient
- |
  patiently
- |
  patina
- |
  patinated
- |
  patination
- |
  patio
- |
  patisserie
- |
  patly
- |
  Patmos
- |
  Patna
- |
  patness
- |
  patois
- |
  Paton
- |
  patriarch
- |
  patriarchal
- |
  patriarchate
- |
  patriarchic
- |
  patriarchy
- |
  patriate
- |
  Patricia
- |
  patrician
- |
  patricidal
- |
  patricide
- |
  Patrick
- |
  patrilineal
- |
  patrimonial
- |
  patrimony
- |
  patriot
- |
  patriotic
- |
  patriotism
- |
  patristic
- |
  patristical
- |
  patrol
- |
  patrolman
- |
  patrolwoman
- |
  patron
- |
  patronage
- |
  patroness
- |
  patronise
- |
  patronising
- |
  patronize
- |
  patronizer
- |
  patronizing
- |
  patronymic
- |
  patroon
- |
  patroonship
- |
  Patsy
- |
  patsy
- |
  patter
- |
  pattern
- |
  patterned
- |
  Patti
- |
  Pattie
- |
  pattie
- |
  Patton
- |
  Patty
- |
  patty
- |
  patulous
- |
  patulously
- |
  patulousness
- |
  paucity
- |
  Paula
- |
  Paulette
- |
  Pauline
- |
  Pauling
- |
  paunch
- |
  paunchy
- |
  pauper
- |
  pauperism
- |
  pauperize
- |
  pause
- |
  pavan
- |
  pavane
- |
  Pavarotti
- |
  paved
- |
  pavement
- |
  pavilion
- |
  paving
- |
  Pavlov
- |
  Pavlova
- |
  Pavlovian
- |
  pawnbroker
- |
  pawnbroking
- |
  Pawnee
- |
  pawnshop
- |
  pawpaw
- |
  payable
- |
  payback
- |
  paycheck
- |
  payday
- |
  payee
- |
  payer
- |
  payload
- |
  paymaster
- |
  payment
- |
  paymistress
- |
  payoff
- |
  payola
- |
  payout
- |
  payroll
- |
  payslip
- |
  peace
- |
  peaceable
- |
  peaceably
- |
  peaceful
- |
  peacefully
- |
  peacefulness
- |
  peacekeeper
- |
  peacekeeping
- |
  peacemaker
- |
  peacemaking
- |
  peacetime
- |
  peach
- |
  peachy
- |
  peacock
- |
  peafowl
- |
  peahen
- |
  peaked
- |
  Peale
- |
  peanut
- |
  peanuts
- |
  Pearl
- |
  pearl
- |
  pearly
- |
  Pearson
- |
  Peary
- |
  peasant
- |
  peasantry
- |
  peashooter
- |
  peatbog
- |
  peatmoss
- |
  peaty
- |
  pebble
- |
  pebbly
- |
  pecan
- |
  peccadillo
- |
  peccancy
- |
  peccant
- |
  peccary
- |
  peccavi
- |
  peckish
- |
  Pecos
- |
  pectic
- |
  pectin
- |
  pectinous
- |
  pectoral
- |
  pectorals
- |
  peculate
- |
  peculation
- |
  peculator
- |
  peculiar
- |
  peculiarity
- |
  peculiarly
- |
  pecuniarily
- |
  pecuniary
- |
  pedagog
- |
  pedagogic
- |
  pedagogical
- |
  pedagogics
- |
  pedagogue
- |
  pedagogy
- |
  pedal
- |
  pedant
- |
  pedantic
- |
  pedantically
- |
  pedantry
- |
  peddle
- |
  peddler
- |
  peddling
- |
  pederast
- |
  pederastic
- |
  pederasty
- |
  pedestal
- |
  pedestrian
- |
  pedestrianly
- |
  pediatric
- |
  pediatrician
- |
  pediatrics
- |
  pedicab
- |
  pedicular
- |
  pediculosis
- |
  pediculous
- |
  pedicure
- |
  pedicurist
- |
  pedigree
- |
  pedigreed
- |
  pediment
- |
  pedimental
- |
  pedimented
- |
  pedlar
- |
  pedological
- |
  pedologist
- |
  pedology
- |
  pedometer
- |
  pedophile
- |
  pedophilia
- |
  pedophilic
- |
  Pedro
- |
  peduncle
- |
  peduncular
- |
  peekaboo
- |
  peeler
- |
  peeling
- |
  peelings
- |
  peeper
- |
  peephole
- |
  peerage
- |
  peeress
- |
  peerless
- |
  peerlessly
- |
  peeve
- |
  peevish
- |
  peevishly
- |
  peevishness
- |
  peewee
- |
  Pegasus
- |
  pegboard
- |
  Peggy
- |
  pegmatite
- |
  peignoir
- |
  Peiping
- |
  pejoration
- |
  pejorative
- |
  pejoratively
- |
  Pekinese
- |
  pekinese
- |
  Peking
- |
  Pekingese
- |
  pekingese
- |
  pekoe
- |
  pelage
- |
  pelagian
- |
  pelagic
- |
  Pelee
- |
  pelican
- |
  Pelion
- |
  pellagra
- |
  pellagrous
- |
  pellet
- |
  pelletal
- |
  pelletize
- |
  pellucid
- |
  pellucidity
- |
  pellucidly
- |
  pellucidness
- |
  Peloponnesus
- |
  Peloponnisos
- |
  pelves
- |
  pelvic
- |
  pelvis
- |
  pemican
- |
  pemmican
- |
  penal
- |
  penalise
- |
  penalization
- |
  penalize
- |
  penally
- |
  penalty
- |
  penance
- |
  Penang
- |
  Penates
- |
  penates
- |
  pence
- |
  penchant
- |
  pencil
- |
  pencilled
- |
  pendant
- |
  pendency
- |
  pendent
- |
  pending
- |
  pendular
- |
  pendulous
- |
  pendulously
- |
  pendulum
- |
  Penelope
- |
  peneplain
- |
  peneplane
- |
  penes
- |
  penetrable
- |
  penetralia
- |
  penetrant
- |
  penetrate
- |
  penetrating
- |
  penetration
- |
  penetrative
- |
  penguin
- |
  penicillin
- |
  penile
- |
  peninsula
- |
  peninsular
- |
  penis
- |
  penitence
- |
  penitent
- |
  penitential
- |
  penitentiary
- |
  penitently
- |
  penknife
- |
  penknives
- |
  penlight
- |
  penlite
- |
  penman
- |
  penmanship
- |
  penname
- |
  pennant
- |
  penne
- |
  penni
- |
  penniless
- |
  Pennines
- |
  pennon
- |
  pennoned
- |
  Pennsylvania
- |
  Penny
- |
  penny
- |
  pennyroyal
- |
  pennyweight
- |
  Penobscot
- |
  penological
- |
  penologist
- |
  penology
- |
  Pensacola
- |
  pensee
- |
  pensile
- |
  pension
- |
  pensionable
- |
  pensioner
- |
  pensive
- |
  pensively
- |
  pensiveness
- |
  penstock
- |
  pentacle
- |
  Pentagon
- |
  pentagon
- |
  pentagonal
- |
  pentagram
- |
  pentameter
- |
  pentangle
- |
  Pentateuch
- |
  Pentateuchal
- |
  pentathlete
- |
  pentathlon
- |
  Pentecost
- |
  Pentecostal
- |
  penthouse
- |
  penuche
- |
  penuchi
- |
  penultimate
- |
  penumbra
- |
  penumbrae
- |
  penumbral
- |
  penurious
- |
  penuriously
- |
  penury
- |
  Penutian
- |
  Penza
- |
  peonage
- |
  peony
- |
  people
- |
  Peoria
- |
  Pepin
- |
  pepper
- |
  peppercorn
- |
  peppermint
- |
  pepperoni
- |
  peppery
- |
  peppiness
- |
  peppy
- |
  pepsin
- |
  peptic
- |
  peptide
- |
  Pepys
- |
  Pepysian
- |
  Pequot
- |
  peradventure
- |
  perambulate
- |
  perambulator
- |
  percale
- |
  perceivable
- |
  perceive
- |
  percent
- |
  percentage
- |
  percentile
- |
  percept
- |
  perceptible
- |
  perceptibly
- |
  perception
- |
  perceptional
- |
  perceptive
- |
  perceptively
- |
  perceptivity
- |
  perceptual
- |
  perceptually
- |
  Perceval
- |
  perch
- |
  perchance
- |
  perched
- |
  percipience
- |
  percipient
- |
  percipiently
- |
  Percival
- |
  percolate
- |
  percolation
- |
  percolator
- |
  percussion
- |
  percussive
- |
  Percy
- |
  perdition
- |
  perdurable
- |
  perdurably
- |
  perdurance
- |
  perdure
- |
  peregrinate
- |
  peregrinator
- |
  peregrine
- |
  peremptorily
- |
  peremptory
- |
  perennial
- |
  perennially
- |
  perestroika
- |
  perfect
- |
  perfecta
- |
  perfectible
- |
  perfection
- |
  perfectly
- |
  perfectness
- |
  perfecto
- |
  perfervid
- |
  perfervidly
- |
  perfidious
- |
  perfidiously
- |
  perfidy
- |
  perforate
- |
  perforated
- |
  perforation
- |
  perforator
- |
  perforce
- |
  perform
- |
  performance
- |
  performative
- |
  performer
- |
  perfume
- |
  perfumed
- |
  perfumer
- |
  perfumery
- |
  perfunctory
- |
  perfuse
- |
  perfusion
- |
  perfusionist
- |
  Pergamum
- |
  Pergamus
- |
  pergola
- |
  perhaps
- |
  perianth
- |
  pericardia
- |
  pericardial
- |
  pericardium
- |
  Periclean
- |
  Pericles
- |
  perigee
- |
  perihelia
- |
  perihelion
- |
  peril
- |
  perilous
- |
  perilously
- |
  perimeter
- |
  perimetric
- |
  perinea
- |
  perineal
- |
  perineum
- |
  period
- |
  periodic
- |
  periodical
- |
  periodically
- |
  periodicity
- |
  periodontal
- |
  periodontics
- |
  periodontist
- |
  Peripatetic
- |
  peripatetic
- |
  peripheral
- |
  peripherally
- |
  periphery
- |
  periphrases
- |
  periphrasis
- |
  periphrastic
- |
  periscope
- |
  periscopic
- |
  perish
- |
  perishable
- |
  perishables
- |
  perishably
- |
  peristalses
- |
  peristalsis
- |
  peristaltic
- |
  peristyle
- |
  peritonea
- |
  peritoneal
- |
  peritoneum
- |
  peritonitis
- |
  periwig
- |
  periwinkle
- |
  perjure
- |
  perjurer
- |
  perjurious
- |
  perjuriously
- |
  perjury
- |
  perkily
- |
  perkiness
- |
  Perkins
- |
  perky
- |
  perlite
- |
  Perlman
- |
  perlocution
- |
  permafrost
- |
  permanence
- |
  permanency
- |
  permanent
- |
  permanently
- |
  permeability
- |
  permeable
- |
  permeate
- |
  permeation
- |
  permeative
- |
  Permian
- |
  permissible
- |
  permissibly
- |
  permission
- |
  permissive
- |
  permissively
- |
  permit
- |
  permitee
- |
  permitter
- |
  permutation
- |
  Pernambuco
- |
  pernicious
- |
  perniciously
- |
  Peron
- |
  perorate
- |
  peroration
- |
  Perot
- |
  peroxide
- |
  perpetrate
- |
  perpetration
- |
  perpetrator
- |
  perpetual
- |
  perpetually
- |
  perpetuance
- |
  perpetuate
- |
  perpetuation
- |
  perpetuator
- |
  perpetuity
- |
  perplex
- |
  perplexed
- |
  perplexedly
- |
  perplexing
- |
  perplexingly
- |
  perplexities
- |
  perplexity
- |
  perquisite
- |
  Perry
- |
  persecute
- |
  persecution
- |
  persecutor
- |
  persecutory
- |
  Persephone
- |
  Persepolis
- |
  Perseus
- |
  perseverance
- |
  perseverate
- |
  persevere
- |
  persevering
- |
  Pershing
- |
  Persia
- |
  Persian
- |
  persiflage
- |
  persimmon
- |
  persist
- |
  persistence
- |
  persistency
- |
  persistent
- |
  persistently
- |
  persnickety
- |
  person
- |
  persona
- |
  personable
- |
  personably
- |
  personae
- |
  personage
- |
  personal
- |
  personalise
- |
  personality
- |
  personalize
- |
  personalized
- |
  personally
- |
  personals
- |
  personalty
- |
  personate
- |
  personifier
- |
  personify
- |
  personnel
- |
  perspective
- |
  perspicacity
- |
  perspicuity
- |
  perspicuous
- |
  perspiration
- |
  perspire
- |
  persuadable
- |
  persuade
- |
  persuaded
- |
  persuader
- |
  persuasible
- |
  persuasion
- |
  persuasive
- |
  persuasively
- |
  pertain
- |
  Perth
- |
  pertinacious
- |
  pertinacity
- |
  pertinence
- |
  pertinency
- |
  pertinent
- |
  pertinently
- |
  pertly
- |
  pertness
- |
  perturb
- |
  perturbable
- |
  perturbation
- |
  perturbative
- |
  perturbed
- |
  perturbingly
- |
  pertussal
- |
  pertussis
- |
  peruke
- |
  perusal
- |
  peruse
- |
  peruser
- |
  Peruvian
- |
  pervade
- |
  pervasion
- |
  pervasive
- |
  pervasively
- |
  perverse
- |
  perversely
- |
  perverseness
- |
  perversion
- |
  perversity
- |
  pervert
- |
  perverted
- |
  perverter
- |
  pervious
- |
  perviously
- |
  perviousness
- |
  peseta
- |
  pesewa
- |
  Peshawar
- |
  peskily
- |
  peskiness
- |
  pesky
- |
  pessimism
- |
  pessimist
- |
  pessimistic
- |
  pester
- |
  pesterer
- |
  pesthole
- |
  pesticide
- |
  pestiferous
- |
  pestilence
- |
  pestilent
- |
  pestilential
- |
  pestle
- |
  pesto
- |
  pesty
- |
  Petain
- |
  petal
- |
  petaled
- |
  petalled
- |
  petard
- |
  petcock
- |
  Peter
- |
  peter
- |
  Peterborough
- |
  petiole
- |
  petit
- |
  petite
- |
  petition
- |
  petitionary
- |
  petitioner
- |
  Petra
- |
  Petrarch
- |
  Petrarchan
- |
  petrel
- |
  petrifaction
- |
  petrified
- |
  petrify
- |
  petrodollar
- |
  petrodollars
- |
  petroglyph
- |
  petroglyphic
- |
  Petrograd
- |
  petrographer
- |
  petrography
- |
  petrol
- |
  petrolatum
- |
  petroleum
- |
  petrologist
- |
  petrology
- |
  petter
- |
  petticoat
- |
  pettifog
- |
  pettifogger
- |
  pettifoggery
- |
  pettily
- |
  pettiness
- |
  pettish
- |
  pettishly
- |
  petty
- |
  petulance
- |
  petulancy
- |
  petulant
- |
  petulantly
- |
  petunia
- |
  pewee
- |
  pewter
- |
  pewterer
- |
  peyote
- |
  peyotl
- |
  pfennig
- |
  pfennige
- |
  phaeton
- |
  phage
- |
  phagocyte
- |
  phagocytic
- |
  phalanger
- |
  phalanges
- |
  phalanx
- |
  phalarope
- |
  phalli
- |
  phallic
- |
  phallically
- |
  phallicism
- |
  phallism
- |
  phallus
- |
  Phanerozoic
- |
  phantasm
- |
  phantasmal
- |
  phantasmic
- |
  phantasy
- |
  phantom
- |
  Pharaoh
- |
  pharaoh
- |
  Pharaonic
- |
  Pharisaic
- |
  pharisaic
- |
  Pharisaical
- |
  pharisaical
- |
  Pharisaism
- |
  Pharisee
- |
  pharisee
- |
  pharmaceutic
- |
  pharmacist
- |
  pharmacology
- |
  pharmacopeia
- |
  pharmacy
- |
  Pharos
- |
  pharos
- |
  pharyngeal
- |
  pharynges
- |
  pharyngitis
- |
  pharyngology
- |
  pharynx
- |
  phase
- |
  phaseout
- |
  phasic
- |
  pheasant
- |
  Phebe
- |
  Phecda
- |
  phenacetin
- |
  phenix
- |
  phenol
- |
  phenolic
- |
  phenom
- |
  phenomena
- |
  phenomenal
- |
  phenomenally
- |
  phenomenon
- |
  phenotype
- |
  phenotypic
- |
  phenotypical
- |
  pheromonal
- |
  pheromone
- |
  phial
- |
  Phidias
- |
  Philadelphia
- |
  philander
- |
  philanderer
- |
  philandering
- |
  philanthropy
- |
  philatelic
- |
  philatelist
- |
  philately
- |
  Philemon
- |
  philharmonic
- |
  Philip
- |
  Philippa
- |
  Philippi
- |
  Philippian
- |
  Philippians
- |
  philippic
- |
  Philippine
- |
  Philippines
- |
  Philistine
- |
  philistine
- |
  philistinish
- |
  philistinism
- |
  Phillip
- |
  Phillips
- |
  Phillis
- |
  philodendra
- |
  philodendron
- |
  philogynist
- |
  philogyny
- |
  philologian
- |
  philological
- |
  philologist
- |
  philology
- |
  philosopher
- |
  philosophic
- |
  philosophize
- |
  philosophy
- |
  philter
- |
  philtre
- |
  Phineas
- |
  phlebitic
- |
  phlebitis
- |
  phlebotomy
- |
  phlegm
- |
  phlegmatic
- |
  phlegmatical
- |
  phlegmy
- |
  phloem
- |
  phlogiston
- |
  phlox
- |
  phobia
- |
  phobic
- |
  Phoebe
- |
  phoebe
- |
  Phoenicia
- |
  Phoenician
- |
  Phoenix
- |
  phoenix
- |
  phone
- |
  phoneme
- |
  phonemic
- |
  phonemically
- |
  phonemics
- |
  phonetic
- |
  phonetically
- |
  phonetician
- |
  phonetics
- |
  phoney
- |
  phonic
- |
  phonically
- |
  phonics
- |
  phoniness
- |
  phonograph
- |
  phonographic
- |
  phonologic
- |
  phonological
- |
  phonologist
- |
  phonology
- |
  phony
- |
  phooey
- |
  phosgene
- |
  phosphate
- |
  phosphatic
- |
  phospholipid
- |
  phosphor
- |
  phosphoresce
- |
  phosphoric
- |
  phosphorous
- |
  phosphorus
- |
  photic
- |
  photo
- |
  photoaging
- |
  photocell
- |
  photocompose
- |
  photocopier
- |
  photocopy
- |
  photoengrave
- |
  photoflash
- |
  photog
- |
  photogenic
- |
  photograph
- |
  photographer
- |
  photographic
- |
  photography
- |
  photogravure
- |
  photometer
- |
  photometric
- |
  photometry
- |
  photomontage
- |
  photon
- |
  photonic
- |
  photoplay
- |
  photorealism
- |
  photorealist
- |
  photosphere
- |
  photospheric
- |
  Photostat
- |
  photostatic
- |
  phototropic
- |
  phototropism
- |
  photovoltaic
- |
  phrasal
- |
  phrase
- |
  phraseology
- |
  phrasing
- |
  phrenetic
- |
  phrenetical
- |
  phrenic
- |
  phrenologic
- |
  phrenologist
- |
  phrenology
- |
  Phrygia
- |
  Phrygian
- |
  phyla
- |
  phylactery
- |
  Phyllis
- |
  phyllo
- |
  phyllotaxes
- |
  phyllotaxis
- |
  phyllotaxy
- |
  phylogenetic
- |
  phylogenic
- |
  phylogenist
- |
  phylogeny
- |
  phylum
- |
  physic
- |
  physical
- |
  physicality
- |
  physically
- |
  physician
- |
  physicist
- |
  physics
- |
  physiognomic
- |
  physiognomy
- |
  physiography
- |
  physiologic
- |
  physiologist
- |
  physiology
- |
  physiotype
- |
  physique
- |
  physiqued
- |
  Piaget
- |
  pianissimi
- |
  pianissimo
- |
  pianist
- |
  piano
- |
  pianoforte
- |
  piaster
- |
  piastre
- |
  piazza
- |
  piazze
- |
  pibroch
- |
  picador
- |
  Picardy
- |
  picaresque
- |
  Picasso
- |
  picayune
- |
  piccalilli
- |
  piccolo
- |
  pickaback
- |
  pickax
- |
  pickaxe
- |
  picked
- |
  picker
- |
  pickerel
- |
  pickerelweed
- |
  picket
- |
  picketer
- |
  picketing
- |
  Pickett
- |
  picking
- |
  pickings
- |
  pickle
- |
  pickled
- |
  pickling
- |
  picklock
- |
  pickpocket
- |
  pickup
- |
  Pickwick
- |
  picky
- |
  picnic
- |
  picnicker
- |
  picot
- |
  pictograph
- |
  pictographic
- |
  Pictor
- |
  pictorial
- |
  pictorially
- |
  picture
- |
  picturesque
- |
  piddle
- |
  piddling
- |
  piddly
- |
  pidgin
- |
  piebald
- |
  piece
- |
  piecemeal
- |
  piecework
- |
  pieceworker
- |
  Piedmont
- |
  piedmont
- |
  Piedmontese
- |
  Pierce
- |
  pierce
- |
  piercing
- |
  piercingly
- |
  Pierre
- |
  Pieta
- |
  pieta
- |
  Pietism
- |
  pietism
- |
  pietist
- |
  pietistic
- |
  pietistical
- |
  piety
- |
  piffle
- |
  piffling
- |
  pigeon
- |
  pigeonhole
- |
  piggish
- |
  piggishly
- |
  piggishness
- |
  piggy
- |
  piggyback
- |
  pigheaded
- |
  piglet
- |
  pigment
- |
  pigmentary
- |
  pigmentation
- |
  Pigmy
- |
  pigmy
- |
  pignut
- |
  pigpen
- |
  pigskin
- |
  pigsty
- |
  pigtail
- |
  pigtailed
- |
  piked
- |
  piker
- |
  pikestaff
- |
  pilaf
- |
  pilaff
- |
  pilaster
- |
  pilastered
- |
  Pilate
- |
  pilau
- |
  pilchard
- |
  piled
- |
  pileless
- |
  piles
- |
  pileup
- |
  pilfer
- |
  pilferage
- |
  pilferer
- |
  Pilgrim
- |
  pilgrim
- |
  pilgrimage
- |
  pilgrimize
- |
  piling
- |
  Pilipino
- |
  pillage
- |
  pillager
- |
  pillaging
- |
  pillar
- |
  pillared
- |
  pillbox
- |
  pillion
- |
  pillory
- |
  pillow
- |
  pillowcase
- |
  pillowslip
- |
  pillowy
- |
  pilose
- |
  pilosity
- |
  pilot
- |
  pilotage
- |
  pilothouse
- |
  pilotless
- |
  pilous
- |
  pilsener
- |
  pilsner
- |
  Piman
- |
  pimento
- |
  pimiento
- |
  pimpernel
- |
  pimping
- |
  pimple
- |
  pimpled
- |
  pimply
- |
  pinafore
- |
  pinata
- |
  pinball
- |
  pincer
- |
  pincers
- |
  pinch
- |
  pinched
- |
  pincher
- |
  pinchers
- |
  pincushion
- |
  Pindar
- |
  Pindaric
- |
  Pindus
- |
  pineal
- |
  pineapple
- |
  piney
- |
  pinfeather
- |
  pinhead
- |
  pinheaded
- |
  pinhole
- |
  pinion
- |
  Pinkerton
- |
  pinkeye
- |
  pinkie
- |
  pinkish
- |
  pinkness
- |
  pinky
- |
  pinnace
- |
  pinnacle
- |
  pinnacled
- |
  pinnate
- |
  pinnated
- |
  pinnately
- |
  pinnation
- |
  Pinocchio
- |
  pinochle
- |
  pinocle
- |
  pinon
- |
  pinones
- |
  pinpoint
- |
  pinprick
- |
  pinsetter
- |
  pinspotter
- |
  pinstripe
- |
  pinstriped
- |
  Pinter
- |
  Pinteresque
- |
  pinto
- |
  pintsize
- |
  pintsized
- |
  pinup
- |
  pinwheel
- |
  pinworm
- |
  Pinyin
- |
  pinyin
- |
  pinyon
- |
  pioneer
- |
  pioneering
- |
  piosity
- |
  pious
- |
  piously
- |
  piousness
- |
  pipeful
- |
  pipeline
- |
  piper
- |
  pipes
- |
  pipestone
- |
  pipet
- |
  pipette
- |
  piping
- |
  pipit
- |
  pippin
- |
  pipsqueak
- |
  piquancy
- |
  piquant
- |
  piquante
- |
  piquantly
- |
  piquantness
- |
  pique
- |
  piquet
- |
  piracy
- |
  Piraeus
- |
  pirana
- |
  Pirandello
- |
  piranha
- |
  pirate
- |
  pirated
- |
  piratic
- |
  piratical
- |
  pirogi
- |
  pirogue
- |
  piroshki
- |
  pirouette
- |
  Pisan
- |
  piscatorial
- |
  piscatory
- |
  Pisces
- |
  pisciculture
- |
  piscina
- |
  piscinae
- |
  piscine
- |
  Pisistratus
- |
  pismire
- |
  Pissaro
- |
  pissed
- |
  pistachio
- |
  pistil
- |
  pistillate
- |
  pistol
- |
  piston
- |
  pitapat
- |
  Pitcairn
- |
  pitch
- |
  pitchblende
- |
  pitcher
- |
  pitcherful
- |
  pitchfork
- |
  pitching
- |
  pitchman
- |
  pitchy
- |
  piteous
- |
  piteously
- |
  piteousness
- |
  pitfall
- |
  pithily
- |
  pithiness
- |
  pithless
- |
  pithy
- |
  pitiable
- |
  pitiableness
- |
  pitiably
- |
  pitiful
- |
  pitifully
- |
  pitifulness
- |
  pitiless
- |
  pitilessly
- |
  pitilessness
- |
  pitman
- |
  piton
- |
  pittance
- |
  pitted
- |
  Pittsburgh
- |
  pituitary
- |
  Piura
- |
  pivot
- |
  pivotal
- |
  pivotally
- |
  pixel
- |
  pixelate
- |
  pixelation
- |
  pixellate
- |
  pixie
- |
  pixilate
- |
  pixilated
- |
  pixilation
- |
  pixillated
- |
  pixyish
- |
  Pizarro
- |
  pizazz
- |
  pizza
- |
  pizzaz
- |
  pizzazz
- |
  pizzeria
- |
  pizzicato
- |
  placable
- |
  placard
- |
  placate
- |
  placater
- |
  placatingly
- |
  placation
- |
  placatory
- |
  Place
- |
  place
- |
  placebo
- |
  placeholder
- |
  placekick
- |
  placekicker
- |
  placement
- |
  placename
- |
  placenta
- |
  placentae
- |
  placental
- |
  placer
- |
  placid
- |
  placidity
- |
  placidly
- |
  placidness
- |
  placings
- |
  placket
- |
  plagiarism
- |
  plagiarist
- |
  plagiarize
- |
  plagiarizer
- |
  plagiary
- |
  plague
- |
  plaice
- |
  plaid
- |
  plain
- |
  plainclothes
- |
  plainly
- |
  plainness
- |
  plainsman
- |
  plainsong
- |
  plainspoken
- |
  plaint
- |
  plaintiff
- |
  plaintive
- |
  plaintively
- |
  plait
- |
  planar
- |
  planarity
- |
  Planck
- |
  plane
- |
  planeload
- |
  planer
- |
  planet
- |
  planetaria
- |
  planetarium
- |
  planetary
- |
  planetesimal
- |
  planetoid
- |
  plangency
- |
  plangent
- |
  plangently
- |
  plank
- |
  planking
- |
  plankton
- |
  planktonic
- |
  planner
- |
  planning
- |
  Plano
- |
  plant
- |
  plantable
- |
  plantain
- |
  plantar
- |
  plantation
- |
  planter
- |
  plantigrade
- |
  planting
- |
  plantlike
- |
  plaque
- |
  plash
- |
  plasm
- |
  plasma
- |
  plasmatic
- |
  plasmic
- |
  plasmin
- |
  plasmolyses
- |
  plasmolysis
- |
  plasmolytic
- |
  plaster
- |
  plasterboard
- |
  plastered
- |
  plasterer
- |
  plastic
- |
  plastically
- |
  plasticity
- |
  plasticize
- |
  plasticizer
- |
  plastid
- |
  plastique
- |
  Plata
- |
  plate
- |
  plateau
- |
  plateaux
- |
  plated
- |
  plateful
- |
  platelet
- |
  platen
- |
  platform
- |
  Plath
- |
  plating
- |
  platinum
- |
  platitude
- |
  Plato
- |
  Platonic
- |
  platonic
- |
  Platonically
- |
  platonically
- |
  Platonism
- |
  Platonist
- |
  platoon
- |
  Platte
- |
  platter
- |
  platy
- |
  platyfish
- |
  platypi
- |
  platypus
- |
  platys
- |
  plaudit
- |
  plaudits
- |
  plausibility
- |
  plausible
- |
  plausibly
- |
  Plautus
- |
  playa
- |
  playable
- |
  playact
- |
  playacting
- |
  playback
- |
  playbill
- |
  playbook
- |
  playboy
- |
  player
- |
  playful
- |
  playfully
- |
  playfulness
- |
  playgirl
- |
  playgoer
- |
  playgoing
- |
  playground
- |
  playgroup
- |
  playhouse
- |
  playlet
- |
  playmate
- |
  playoff
- |
  playpen
- |
  playroom
- |
  playsuit
- |
  plaything
- |
  playwright
- |
  plaza
- |
  plead
- |
  pleader
- |
  pleading
- |
  pleadingly
- |
  pleasant
- |
  pleasantly
- |
  pleasantness
- |
  pleasantry
- |
  please
- |
  pleased
- |
  pleasing
- |
  pleasingly
- |
  pleasurable
- |
  pleasurably
- |
  pleasure
- |
  pleasureful
- |
  pleat
- |
  pleated
- |
  plebe
- |
  plebeian
- |
  plebes
- |
  plebiscitary
- |
  plebiscite
- |
  plebs
- |
  plectra
- |
  plectrum
- |
  pledge
- |
  pledger
- |
  pleiad
- |
  Pleiades
- |
  Pleistocene
- |
  plena
- |
  plenarily
- |
  plenary
- |
  plenitude
- |
  plenteous
- |
  plentiful
- |
  plentifully
- |
  plenty
- |
  plenum
- |
  pleonasm
- |
  pleonastic
- |
  plesiosaur
- |
  plesiosaurus
- |
  plethora
- |
  plethoric
- |
  pleura
- |
  pleurae
- |
  pleural
- |
  pleurisy
- |
  pleuritic
- |
  plexiform
- |
  Plexiglas
- |
  Plexiglass
- |
  plexiglass
- |
  plexus
- |
  pliability
- |
  pliable
- |
  pliableness
- |
  pliably
- |
  pliancy
- |
  pliant
- |
  pliers
- |
  plight
- |
  plighter
- |
  plinth
- |
  Pliny
- |
  Pliocene
- |
  plodder
- |
  plodding
- |
  ploddingly
- |
  Ploesti
- |
  plosion
- |
  plosive
- |
  plotter
- |
  plough
- |
  ploughing
- |
  Plovdiv
- |
  plover
- |
  plowable
- |
  plowboy
- |
  plower
- |
  plowing
- |
  plowman
- |
  plowshare
- |
  pluck
- |
  pluckily
- |
  pluckiness
- |
  plucky
- |
  plugola
- |
  plumage
- |
  plumaged
- |
  plumb
- |
  plumbable
- |
  plumber
- |
  plumbing
- |
  plume
- |
  plumed
- |
  plummet
- |
  plummy
- |
  plump
- |
  plumpness
- |
  plumy
- |
  plunder
- |
  plunderer
- |
  plunge
- |
  plunger
- |
  plunk
- |
  plunker
- |
  pluperfect
- |
  plural
- |
  pluralism
- |
  pluralist
- |
  pluralistic
- |
  plurality
- |
  pluralize
- |
  plush
- |
  plushily
- |
  plushiness
- |
  plushly
- |
  plushness
- |
  plushy
- |
  Plutarch
- |
  Pluto
- |
  plutocracy
- |
  plutocrat
- |
  plutocratic
- |
  plutonic
- |
  plutonium
- |
  pluvial
- |
  Plymouth
- |
  plywood
- |
  pneumatic
- |
  pneumatical
- |
  pneumaticity
- |
  pneumatics
- |
  pneumococcal
- |
  pneumococci
- |
  pneumococcus
- |
  pneumonia
- |
  pneumonic
- |
  poach
- |
  poacher
- |
  Pocahontas
- |
  Pocatello
- |
  pocked
- |
  pocket
- |
  pocketbook
- |
  pocketful
- |
  pocketknife
- |
  pocketknives
- |
  pockmark
- |
  pockmarked
- |
  Podgorica
- |
  podia
- |
  podiatric
- |
  podiatrist
- |
  podiatry
- |
  podium
- |
  poesy
- |
  poetaster
- |
  poetess
- |
  poetic
- |
  poetical
- |
  poetically
- |
  poetry
- |
  pogrom
- |
  poignance
- |
  poignancy
- |
  poignant
- |
  poignantly
- |
  poikilotherm
- |
  poinciana
- |
  poinsettia
- |
  point
- |
  pointed
- |
  pointedly
- |
  pointelle
- |
  pointer
- |
  pointillism
- |
  pointillist
- |
  pointilliste
- |
  pointless
- |
  pointlessly
- |
  pointy
- |
  poise
- |
  poised
- |
  poisha
- |
  poison
- |
  poisoned
- |
  poisoner
- |
  poisoning
- |
  poisonous
- |
  poisonously
- |
  poker
- |
  pokeweed
- |
  pokey
- |
  pokily
- |
  pokiness
- |
  Poland
- |
  polar
- |
  Polaris
- |
  polarise
- |
  polarity
- |
  polarizable
- |
  polarization
- |
  polarize
- |
  polarized
- |
  polarizer
- |
  polarizing
- |
  Polaroid
- |
  polder
- |
  poleax
- |
  poleaxe
- |
  polecat
- |
  polemic
- |
  polemical
- |
  polemicist
- |
  polemicize
- |
  polemics
- |
  polenta
- |
  poler
- |
  polestar
- |
  poleward
- |
  police
- |
  policeman
- |
  policewoman
- |
  policing
- |
  policy
- |
  policyholder
- |
  policymaker
- |
  policymaking
- |
  polio
- |
  Polish
- |
  polish
- |
  polished
- |
  polisher
- |
  Politburo
- |
  politburo
- |
  polite
- |
  politely
- |
  politeness
- |
  politesse
- |
  politic
- |
  political
- |
  politically
- |
  politician
- |
  politicise
- |
  politicize
- |
  politicized
- |
  politick
- |
  politicker
- |
  politicking
- |
  politicly
- |
  politico
- |
  politics
- |
  polity
- |
  polka
- |
  pollack
- |
  pollen
- |
  poller
- |
  pollinate
- |
  pollination
- |
  pollinator
- |
  polling
- |
  pollinosis
- |
  polliwog
- |
  Pollock
- |
  pollock
- |
  polls
- |
  pollster
- |
  pollutant
- |
  pollute
- |
  polluted
- |
  polluter
- |
  pollution
- |
  Pollux
- |
  Polly
- |
  Pollyanna
- |
  pollywog
- |
  polonaise
- |
  polonium
- |
  poltergeist
- |
  poltroon
- |
  poltroonery
- |
  poltroonish
- |
  polyandrous
- |
  polyandry
- |
  polychrome
- |
  polychromed
- |
  polychromic
- |
  polychromous
- |
  polyclinic
- |
  polydipsia
- |
  polydipsic
- |
  polyester
- |
  polyethylene
- |
  polygamist
- |
  polygamous
- |
  polygamously
- |
  polygamy
- |
  polyglot
- |
  polyglotism
- |
  polygon
- |
  polygonal
- |
  polygraph
- |
  polygrapher
- |
  polygraphic
- |
  polygynous
- |
  polygyny
- |
  polyhedra
- |
  polyhedral
- |
  polyhedron
- |
  polymath
- |
  polymathic
- |
  polymathy
- |
  polymer
- |
  polymerase
- |
  polymeric
- |
  polymerize
- |
  Polynesia
- |
  Polynesian
- |
  polynomial
- |
  polyp
- |
  polypeptide
- |
  Polyphemus
- |
  polyphonic
- |
  polyphonous
- |
  polyphony
- |
  polypoid
- |
  polys
- |
  polystyrene
- |
  polysyllabic
- |
  polysyllable
- |
  polytechnic
- |
  polytheism
- |
  polytheist
- |
  polytheistic
- |
  polythene
- |
  polyurethane
- |
  polyvalence
- |
  polyvalency
- |
  polyvalent
- |
  polyvinyl
- |
  pomade
- |
  pomander
- |
  pomegranate
- |
  Pomerania
- |
  Pomeranian
- |
  pommel
- |
  Pomona
- |
  Pompadour
- |
  pompadour
- |
  pompano
- |
  Pompeian
- |
  Pompeii
- |
  Pompeiian
- |
  Pompey
- |
  Pompidou
- |
  pompom
- |
  pompon
- |
  pomposity
- |
  pompous
- |
  pompously
- |
  pompousness
- |
  Ponape
- |
  Ponce
- |
  poncho
- |
  ponder
- |
  ponderable
- |
  ponderer
- |
  ponderosa
- |
  ponderosity
- |
  ponderous
- |
  ponderously
- |
  Pondicherry
- |
  Pondoland
- |
  pongee
- |
  poniard
- |
  pontes
- |
  Pontiac
- |
  Pontianak
- |
  Pontic
- |
  pontiff
- |
  pontifical
- |
  pontifically
- |
  pontificals
- |
  Pontificate
- |
  pontificate
- |
  pontificator
- |
  pontoon
- |
  Pontus
- |
  ponytail
- |
  pooch
- |
  poodle
- |
  Poole
- |
  poolroom
- |
  Poona
- |
  pooped
- |
  poorhouse
- |
  poorly
- |
  poormouth
- |
  poorness
- |
  popcorn
- |
  popeyed
- |
  popgun
- |
  popinjay
- |
  poplar
- |
  poplin
- |
  Popocatepetl
- |
  popover
- |
  poppa
- |
  popper
- |
  poppy
- |
  poppycock
- |
  Popsicle
- |
  populace
- |
  popular
- |
  popularise
- |
  popularity
- |
  popularize
- |
  popularizer
- |
  popularly
- |
  populate
- |
  populated
- |
  population
- |
  populism
- |
  populist
- |
  populistic
- |
  populous
- |
  populousness
- |
  porcelain
- |
  porch
- |
  porcine
- |
  porcupine
- |
  pored
- |
  porker
- |
  porky
- |
  porno
- |
  pornographer
- |
  pornographic
- |
  pornography
- |
  porosity
- |
  porous
- |
  porously
- |
  porousness
- |
  porphyritic
- |
  porphyry
- |
  porpoise
- |
  porridge
- |
  porringer
- |
  Porsche
- |
  portability
- |
  portable
- |
  portableness
- |
  portably
- |
  portage
- |
  portal
- |
  portaled
- |
  portalled
- |
  portamenti
- |
  portamento
- |
  portcullis
- |
  portend
- |
  portent
- |
  portentous
- |
  portentously
- |
  Porter
- |
  porter
- |
  porterhouse
- |
  portfolio
- |
  porthole
- |
  Portia
- |
  portico
- |
  portiere
- |
  portion
- |
  Portland
- |
  Portlander
- |
  portliness
- |
  portly
- |
  portmanteau
- |
  portmanteaux
- |
  Porto
- |
  portrait
- |
  portraitist
- |
  portraiture
- |
  portray
- |
  portrayal
- |
  portrayer
- |
  Portsmouth
- |
  Portugal
- |
  Portuguese
- |
  portulaca
- |
  posable
- |
  Poseidon
- |
  poser
- |
  poseur
- |
  poshly
- |
  poshness
- |
  posit
- |
  position
- |
  positional
- |
  positioner
- |
  positive
- |
  positively
- |
  positiveness
- |
  positivism
- |
  positivist
- |
  positivistic
- |
  positivity
- |
  positron
- |
  posse
- |
  possess
- |
  possessed
- |
  possession
- |
  possessions
- |
  possessive
- |
  possessively
- |
  possessor
- |
  possibility
- |
  possible
- |
  possibly
- |
  possum
- |
  postage
- |
  postal
- |
  postally
- |
  postcard
- |
  postcoital
- |
  postcolonial
- |
  postdate
- |
  postdoctoral
- |
  postelection
- |
  poster
- |
  posterior
- |
  posteriority
- |
  posteriorly
- |
  posterity
- |
  postern
- |
  postglacial
- |
  postgraduate
- |
  posthaste
- |
  posthole
- |
  posthumous
- |
  posthumously
- |
  posthypnotic
- |
  postilion
- |
  postillion
- |
  posting
- |
  postlaunch
- |
  postlude
- |
  postman
- |
  postmarital
- |
  postmark
- |
  postmaster
- |
  postmeridian
- |
  postmistress
- |
  postmodern
- |
  postmortem
- |
  postnasal
- |
  postnatal
- |
  postnatally
- |
  postnuptial
- |
  postorgasmic
- |
  postpaid
- |
  postpartum
- |
  postponable
- |
  postpone
- |
  postponement
- |
  postponer
- |
  postprandial
- |
  postscript
- |
  postseason
- |
  postseasonal
- |
  postulancy
- |
  postulant
- |
  postulate
- |
  postulation
- |
  postural
- |
  posture
- |
  posturer
- |
  posturing
- |
  posturist
- |
  postwar
- |
  potability
- |
  potable
- |
  potables
- |
  potage
- |
  potash
- |
  potassic
- |
  potassium
- |
  potation
- |
  potato
- |
  Potawatomi
- |
  potbellied
- |
  potbelly
- |
  potboiler
- |
  potence
- |
  potency
- |
  potent
- |
  potentate
- |
  potential
- |
  potentiality
- |
  potentially
- |
  potentiate
- |
  potentiation
- |
  potently
- |
  potful
- |
  pothead
- |
  pother
- |
  potherb
- |
  potholder
- |
  pothole
- |
  potholed
- |
  pothook
- |
  potion
- |
  potluck
- |
  Potomac
- |
  potpie
- |
  potpourri
- |
  Potsdam
- |
  potshard
- |
  potsherd
- |
  potshot
- |
  pottage
- |
  potted
- |
  Potter
- |
  potter
- |
  pottery
- |
  potty
- |
  pouch
- |
  Poughkeepsie
- |
  poult
- |
  poulterer
- |
  poultice
- |
  poultry
- |
  poultryman
- |
  pounce
- |
  pouncer
- |
  Pound
- |
  pound
- |
  poundage
- |
  poundcake
- |
  pounder
- |
  pounding
- |
  pourboire
- |
  pourer
- |
  pouter
- |
  poutingly
- |
  pouty
- |
  poverty
- |
  powder
- |
  powdered
- |
  powdery
- |
  Powell
- |
  power
- |
  powerboat
- |
  powerful
- |
  powerfully
- |
  powerfulness
- |
  powerhouse
- |
  powerless
- |
  powerlessly
- |
  powers
- |
  powertrain
- |
  Powhatan
- |
  powwow
- |
  Powys
- |
  Poznan
- |
  practicable
- |
  practicably
- |
  practical
- |
  practicality
- |
  practically
- |
  practice
- |
  practiced
- |
  practicer
- |
  practicing
- |
  practicum
- |
  practise
- |
  practising
- |
  practitioner
- |
  Prado
- |
  praesidium
- |
  praetor
- |
  Praetorian
- |
  praetorian
- |
  pragmatic
- |
  pragmatical
- |
  pragmatics
- |
  pragmatism
- |
  pragmatist
- |
  pragmatistic
- |
  Prague
- |
  Praia
- |
  prairie
- |
  praise
- |
  praiseworthy
- |
  praline
- |
  prance
- |
  prancer
- |
  prancingly
- |
  prandial
- |
  prank
- |
  prankster
- |
  praseodymium
- |
  prate
- |
  prater
- |
  pratfall
- |
  prattle
- |
  prattler
- |
  prawn
- |
  praxes
- |
  praxis
- |
  Praxiteles
- |
  prayer
- |
  prayerful
- |
  prayerfully
- |
  prayers
- |
  preach
- |
  preacher
- |
  preachment
- |
  preachy
- |
  preadapt
- |
  preaddress
- |
  preadjust
- |
  preadmission
- |
  preadult
- |
  preamble
- |
  preambular
- |
  preambulary
- |
  preamplifier
- |
  preannounce
- |
  preapply
- |
  preappoint
- |
  preapprove
- |
  prearrange
- |
  prearranged
- |
  preassemble
- |
  preassign
- |
  preassigned
- |
  prebake
- |
  prebend
- |
  prebendary
- |
  preboil
- |
  prebook
- |
  prebuilt
- |
  precalculate
- |
  Precambrian
- |
  precancel
- |
  precancerous
- |
  precarious
- |
  precariously
- |
  precatory
- |
  precaution
- |
  precede
- |
  precedence
- |
  precedent
- |
  preceding
- |
  precentor
- |
  precept
- |
  preceptive
- |
  preceptor
- |
  preceptorial
- |
  precess
- |
  precession
- |
  precessional
- |
  prechill
- |
  precinct
- |
  precincts
- |
  preciosity
- |
  precious
- |
  preciously
- |
  preciousness
- |
  precipice
- |
  precipitable
- |
  precipitance
- |
  precipitancy
- |
  precipitant
- |
  precipitate
- |
  precipitator
- |
  precipitous
- |
  precis
- |
  precise
- |
  precisely
- |
  preciseness
- |
  precision
- |
  preclean
- |
  preclude
- |
  preclusion
- |
  preclusive
- |
  preclusively
- |
  precocious
- |
  precociously
- |
  precocity
- |
  precognition
- |
  precognitive
- |
  precollege
- |
  precolonial
- |
  preconceive
- |
  preconceived
- |
  preconcerted
- |
  precondition
- |
  preconscious
- |
  precook
- |
  precool
- |
  precursor
- |
  precursory
- |
  precut
- |
  predaceous
- |
  predacious
- |
  predacity
- |
  predate
- |
  predation
- |
  predator
- |
  predatorily
- |
  predatory
- |
  predawn
- |
  predecease
- |
  predecessor
- |
  predesignate
- |
  predestinate
- |
  predestine
- |
  predestined
- |
  predetermine
- |
  predicable
- |
  predicament
- |
  predicate
- |
  predication
- |
  predicative
- |
  predict
- |
  predictable
- |
  predictably
- |
  prediction
- |
  predictive
- |
  predictor
- |
  predigest
- |
  predigestion
- |
  predilection
- |
  predinner
- |
  predispose
- |
  predisposed
- |
  predominance
- |
  predominancy
- |
  predominant
- |
  predominate
- |
  predominator
- |
  preelection
- |
  preemie
- |
  preeminence
- |
  preeminent
- |
  preeminently
- |
  preempt
- |
  preemption
- |
  preemptive
- |
  preemptor
- |
  preen
- |
  preengage
- |
  preestablish
- |
  preexamine
- |
  preexist
- |
  preexistence
- |
  preexistent
- |
  preexisting
- |
  preexpose
- |
  preexposure
- |
  prefab
- |
  prefabricate
- |
  preface
- |
  prefatory
- |
  prefect
- |
  prefectoral
- |
  prefectorial
- |
  prefectural
- |
  prefecture
- |
  prefer
- |
  preferable
- |
  preferably
- |
  preference
- |
  preferential
- |
  preferment
- |
  prefigure
- |
  prefix
- |
  preflight
- |
  preform
- |
  prefrontal
- |
  pregame
- |
  preglacial
- |
  pregnability
- |
  pregnable
- |
  pregnancy
- |
  pregnant
- |
  pregnantly
- |
  preharden
- |
  preheat
- |
  prehensile
- |
  prehensility
- |
  prehistoric
- |
  prehistory
- |
  prehominid
- |
  prehuman
- |
  preignition
- |
  preinaugural
- |
  preinsert
- |
  preinstruct
- |
  prejudge
- |
  prejudgment
- |
  prejudice
- |
  prejudiced
- |
  prejudicial
- |
  prelacy
- |
  prelate
- |
  prelatic
- |
  prelatical
- |
  prelaunch
- |
  prelim
- |
  preliminary
- |
  preliterate
- |
  prelude
- |
  preludial
- |
  premarital
- |
  premature
- |
  prematurely
- |
  premed
- |
  premedical
- |
  premeditate
- |
  premeditated
- |
  premenstrual
- |
  premie
- |
  Premier
- |
  premier
- |
  premiere
- |
  premiership
- |
  premigration
- |
  premise
- |
  premises
- |
  premium
- |
  premix
- |
  premodern
- |
  premolar
- |
  premonition
- |
  premonitory
- |
  prenatal
- |
  prenatally
- |
  prenotify
- |
  prenuptial
- |
  preoccupied
- |
  preoccupy
- |
  preoperative
- |
  preordain
- |
  preordained
- |
  preowned
- |
  prepackage
- |
  prepaid
- |
  preparation
- |
  preparations
- |
  preparatory
- |
  prepare
- |
  prepared
- |
  preparedness
- |
  prepay
- |
  prepayment
- |
  preplan
- |
  preponderant
- |
  preponderate
- |
  preposition
- |
  prepossess
- |
  preposterous
- |
  preppie
- |
  preppiness
- |
  preppy
- |
  preprandial
- |
  preprogram
- |
  prepuberty
- |
  prepubescent
- |
  prepuce
- |
  preputial
- |
  prequel
- |
  prerecord
- |
  prerecorded
- |
  preregister
- |
  prerelease
- |
  prerequisite
- |
  prerogative
- |
  presage
- |
  presager
- |
  presbyopia
- |
  presbyopic
- |
  presbyter
- |
  presbyteral
- |
  presbyterate
- |
  presbyterial
- |
  Presbyterian
- |
  presbyterian
- |
  presbytery
- |
  preschool
- |
  preschooler
- |
  prescience
- |
  prescient
- |
  presciently
- |
  prescind
- |
  Prescott
- |
  prescreen
- |
  prescreening
- |
  prescribe
- |
  prescriber
- |
  prescript
- |
  prescription
- |
  prescriptive
- |
  preseason
- |
  preselect
- |
  presence
- |
  present
- |
  presentable
- |
  presentably
- |
  presentation
- |
  presenter
- |
  presentient
- |
  presentiment
- |
  presently
- |
  presentment
- |
  presentness
- |
  presents
- |
  preservable
- |
  preservation
- |
  preservative
- |
  preserve
- |
  preserver
- |
  preserves
- |
  preset
- |
  preshrank
- |
  preshrink
- |
  preshrunk
- |
  preshrunken
- |
  preside
- |
  presidency
- |
  President
- |
  president
- |
  presidential
- |
  presidia
- |
  presidio
- |
  Presidium
- |
  presidium
- |
  presignify
- |
  preslavery
- |
  Presley
- |
  presoak
- |
  presort
- |
  press
- |
  pressed
- |
  presser
- |
  pressing
- |
  pressingly
- |
  pressman
- |
  pressroom
- |
  pressure
- |
  pressured
- |
  pressurised
- |
  pressurize
- |
  pressurized
- |
  pressurizer
- |
  prestige
- |
  prestigeful
- |
  prestigious
- |
  presto
- |
  Preston
- |
  prestress
- |
  presumable
- |
  presumably
- |
  presume
- |
  presumption
- |
  presumptive
- |
  presumptuous
- |
  presuppose
- |
  presurgical
- |
  pretax
- |
  preteen
- |
  pretence
- |
  pretend
- |
  pretender
- |
  pretense
- |
  pretension
- |
  pretensions
- |
  pretentious
- |
  preterit
- |
  preterite
- |
  preterm
- |
  pretest
- |
  pretext
- |
  Pretoria
- |
  pretreat
- |
  pretreatment
- |
  pretrial
- |
  prettify
- |
  prettily
- |
  prettiness
- |
  pretty
- |
  pretzel
- |
  prevail
- |
  prevailer
- |
  prevailing
- |
  prevailingly
- |
  prevalence
- |
  prevalent
- |
  prevalently
- |
  prevaricate
- |
  prevaricator
- |
  prevent
- |
  preventable
- |
  preventative
- |
  preventible
- |
  prevention
- |
  preventive
- |
  preverbal
- |
  preview
- |
  Previn
- |
  previous
- |
  previously
- |
  previousness
- |
  prevision
- |
  prevue
- |
  prewar
- |
  prewarm
- |
  prewash
- |
  prexy
- |
  Priam
- |
  priapean
- |
  priapic
- |
  priapism
- |
  Pribilof
- |
  Price
- |
  price
- |
  priceless
- |
  pricey
- |
  pricing
- |
  prick
- |
  pricker
- |
  prickle
- |
  prickliness
- |
  prickly
- |
  pricy
- |
  pride
- |
  prideful
- |
  pridefully
- |
  pridefulness
- |
  prier
- |
  priest
- |
  priestess
- |
  priesthood
- |
  Priestley
- |
  priestliness
- |
  priestly
- |
  priggery
- |
  priggish
- |
  priggishly
- |
  priggishness
- |
  primacy
- |
  primaeval
- |
  primal
- |
  primally
- |
  primarily
- |
  primary
- |
  primate
- |
  primatial
- |
  prime
- |
  primeness
- |
  primer
- |
  primetime
- |
  primeval
- |
  primevally
- |
  primitive
- |
  primitively
- |
  primitivism
- |
  primitivist
- |
  primitivity
- |
  primly
- |
  primness
- |
  primogenital
- |
  primogenitor
- |
  primordial
- |
  primordially
- |
  primp
- |
  primrose
- |
  prince
- |
  princedom
- |
  princeliness
- |
  princeling
- |
  princely
- |
  princess
- |
  Princeton
- |
  principal
- |
  principality
- |
  principally
- |
  Principe
- |
  principle
- |
  principled
- |
  principles
- |
  prink
- |
  prinker
- |
  print
- |
  printable
- |
  printer
- |
  printhead
- |
  printing
- |
  printmaker
- |
  printmaking
- |
  printout
- |
  printwheel
- |
  prior
- |
  priorate
- |
  prioress
- |
  prioritize
- |
  priority
- |
  priorship
- |
  priory
- |
  Priscilla
- |
  prise
- |
  prism
- |
  prismatic
- |
  prison
- |
  prisoner
- |
  prissily
- |
  prissiness
- |
  prissy
- |
  Pristina
- |
  pristine
- |
  pristinely
- |
  prithee
- |
  privacy
- |
  Private
- |
  private
- |
  privateer
- |
  privateering
- |
  privately
- |
  privateness
- |
  privates
- |
  privation
- |
  privatise
- |
  privatize
- |
  privet
- |
  privilege
- |
  privileged
- |
  privily
- |
  privity
- |
  privy
- |
  prize
- |
  prized
- |
  prizefight
- |
  prizefighter
- |
  prizewinner
- |
  prizewinning
- |
  proabortion
- |
  proaction
- |
  proactive
- |
  proactively
- |
  proactivity
- |
  probabilism
- |
  probability
- |
  probable
- |
  probably
- |
  probate
- |
  probation
- |
  probational
- |
  probationary
- |
  probationer
- |
  probative
- |
  probe
- |
  probing
- |
  probity
- |
  problem
- |
  problematic
- |
  probosces
- |
  proboscides
- |
  proboscis
- |
  probusiness
- |
  procaine
- |
  procaryote
- |
  procedural
- |
  procedurally
- |
  procedure
- |
  proceed
- |
  proceeding
- |
  proceedings
- |
  proceeds
- |
  process
- |
  processing
- |
  procession
- |
  processional
- |
  processor
- |
  prochurch
- |
  proclaim
- |
  proclamation
- |
  proclerical
- |
  proclivity
- |
  procommunism
- |
  procommunist
- |
  proconsul
- |
  proconsular
- |
  procreant
- |
  procreate
- |
  procreation
- |
  procreative
- |
  procreator
- |
  Procrustean
- |
  procrustean
- |
  Procrustes
- |
  proctologist
- |
  proctology
- |
  proctor
- |
  proctorial
- |
  procurable
- |
  procurator
- |
  procure
- |
  procurement
- |
  procurer
- |
  procuress
- |
  Procyon
- |
  prodder
- |
  prodding
- |
  prodigal
- |
  prodigality
- |
  prodigally
- |
  prodigious
- |
  prodigiously
- |
  prodigy
- |
  produce
- |
  producer
- |
  producible
- |
  product
- |
  production
- |
  productive
- |
  productively
- |
  productivity
- |
  proem
- |
  proemial
- |
  profanation
- |
  profanatory
- |
  profane
- |
  profanely
- |
  profaneness
- |
  profaner
- |
  profanity
- |
  profascist
- |
  profeminist
- |
  profess
- |
  professed
- |
  professedly
- |
  profession
- |
  professional
- |
  professor
- |
  professorial
- |
  proffer
- |
  proficiency
- |
  proficient
- |
  proficiently
- |
  profile
- |
  profit
- |
  profitable
- |
  profitably
- |
  profiteer
- |
  profiteering
- |
  profiterole
- |
  profitless
- |
  profits
- |
  profligacy
- |
  profligate
- |
  profligately
- |
  profound
- |
  profoundly
- |
  profoundness
- |
  profundity
- |
  profuse
- |
  profusely
- |
  profuseness
- |
  profusion
- |
  progenitive
- |
  progenitor
- |
  progeny
- |
  progesterone
- |
  prognathism
- |
  prognathous
- |
  prognoses
- |
  prognosis
- |
  prognostic
- |
  program
- |
  programer
- |
  programing
- |
  programmable
- |
  programmatic
- |
  programme
- |
  programmer
- |
  programming
- |
  progress
- |
  progression
- |
  progressive
- |
  progun
- |
  prohibit
- |
  Prohibition
- |
  prohibition
- |
  prohibitive
- |
  prohibitor
- |
  prohibitory
- |
  proindustry
- |
  project
- |
  projectile
- |
  projection
- |
  projector
- |
  prokaryote
- |
  prokaryotic
- |
  Prokofiev
- |
  prolabor
- |
  prolapse
- |
  prolate
- |
  prole
- |
  prolegomena
- |
  prolegomenon
- |
  prolepses
- |
  prolepsis
- |
  proleptic
- |
  proletarian
- |
  proletariat
- |
  proliferate
- |
  proliferator
- |
  prolific
- |
  prolificacy
- |
  prolifically
- |
  prolificness
- |
  prolix
- |
  prolixity
- |
  prolixly
- |
  prolog
- |
  prologue
- |
  prolong
- |
  prolongate
- |
  prolongation
- |
  prolonged
- |
  prolusion
- |
  promenade
- |
  Promethean
- |
  Prometheus
- |
  promethium
- |
  promilitary
- |
  prominence
- |
  prominent
- |
  prominently
- |
  promiscuity
- |
  promiscuous
- |
  promise
- |
  promiser
- |
  promising
- |
  promisingly
- |
  promissory
- |
  promo
- |
  promodern
- |
  Promontory
- |
  promontory
- |
  promote
- |
  promoter
- |
  promotion
- |
  promotional
- |
  prompt
- |
  promptbook
- |
  prompter
- |
  prompting
- |
  promptitude
- |
  promptly
- |
  promptness
- |
  promulgate
- |
  promulgation
- |
  promulgator
- |
  pronate
- |
  pronated
- |
  pronation
- |
  pronator
- |
  prone
- |
  proneness
- |
  prong
- |
  pronged
- |
  pronghorn
- |
  pronominal
- |
  pronoun
- |
  pronounce
- |
  pronounced
- |
  pronouncedly
- |
  pronto
- |
  pronuclear
- |
  proof
- |
  proofread
- |
  proofreader
- |
  propaedeutic
- |
  propaganda
- |
  propagandist
- |
  propagandize
- |
  propagate
- |
  propagation
- |
  propagative
- |
  propagator
- |
  propane
- |
  propel
- |
  propellant
- |
  propellent
- |
  propeller
- |
  propellor
- |
  propensity
- |
  proper
- |
  properly
- |
  properness
- |
  propertied
- |
  property
- |
  prophecy
- |
  prophesier
- |
  prophesy
- |
  Prophet
- |
  prophet
- |
  prophetess
- |
  prophetic
- |
  prophetical
- |
  Prophets
- |
  prophylactic
- |
  prophylaxes
- |
  prophylaxis
- |
  propinquity
- |
  propitiate
- |
  propitiation
- |
  propitiator
- |
  propitiatory
- |
  propitious
- |
  propitiously
- |
  propman
- |
  proponent
- |
  proportion
- |
  proportional
- |
  proportions
- |
  proposal
- |
  propose
- |
  proposer
- |
  proposition
- |
  propound
- |
  propounder
- |
  proprietary
- |
  proprieties
- |
  proprietor
- |
  proprietress
- |
  propriety
- |
  propulsion
- |
  propulsive
- |
  prorate
- |
  proration
- |
  proreform
- |
  prorogation
- |
  prorogue
- |
  prosaic
- |
  prosaically
- |
  prosaicness
- |
  proscenia
- |
  proscenium
- |
  prosciutti
- |
  prosciutto
- |
  proscribe
- |
  proscription
- |
  proscriptive
- |
  prose
- |
  prosecutable
- |
  prosecute
- |
  prosecution
- |
  prosecutor
- |
  proselyte
- |
  proselytism
- |
  proselytize
- |
  proselytizer
- |
  prosimian
- |
  prosiness
- |
  proslavery
- |
  prosodic
- |
  prosodical
- |
  prosodist
- |
  prosody
- |
  prospect
- |
  prospecting
- |
  prospective
- |
  prospector
- |
  prospects
- |
  prospectus
- |
  prosper
- |
  prosperity
- |
  prosperous
- |
  prosperously
- |
  prostate
- |
  prostatic
- |
  prostatitis
- |
  prostheses
- |
  prosthesis
- |
  prosthetic
- |
  prostitute
- |
  prostitution
- |
  prostrate
- |
  prostration
- |
  prosy
- |
  protactinium
- |
  protagonist
- |
  Protagoras
- |
  Protagorean
- |
  protean
- |
  proteanism
- |
  protect
- |
  protected
- |
  protection
- |
  protective
- |
  protectively
- |
  Protector
- |
  protector
- |
  Protectorate
- |
  protectorate
- |
  protege
- |
  protegee
- |
  protein
- |
  Proterozoic
- |
  protest
- |
  Protestant
- |
  protestant
- |
  protestation
- |
  protester
- |
  protestor
- |
  Proteus
- |
  prothalmia
- |
  prothalmion
- |
  prothalmium
- |
  protocol
- |
  proton
- |
  protonic
- |
  protoplasm
- |
  protoplasmic
- |
  prototypal
- |
  prototype
- |
  prototypic
- |
  prototypical
- |
  protozoa
- |
  protozoan
- |
  protozoic
- |
  protozoon
- |
  protract
- |
  protracted
- |
  protractile
- |
  protraction
- |
  protractor
- |
  protrude
- |
  protruding
- |
  protrusile
- |
  protrusion
- |
  protrusive
- |
  protuberance
- |
  protuberant
- |
  proud
- |
  Proudhon
- |
  proudly
- |
  proudness
- |
  Proust
- |
  Proustian
- |
  provability
- |
  provable
- |
  prove
- |
  proven
- |
  provenance
- |
  Provencal
- |
  Provence
- |
  provender
- |
  provenience
- |
  proverb
- |
  proverbial
- |
  proverbially
- |
  Proverbs
- |
  provide
- |
  provided
- |
  Providence
- |
  providence
- |
  provident
- |
  providential
- |
  providently
- |
  provider
- |
  providing
- |
  province
- |
  provinces
- |
  provincial
- |
  provincially
- |
  provision
- |
  provisional
- |
  provisioner
- |
  provisions
- |
  proviso
- |
  provisory
- |
  Provo
- |
  provocation
- |
  provocative
- |
  provoke
- |
  provoker
- |
  provoking
- |
  provolone
- |
  provost
- |
  provostship
- |
  prowess
- |
  prowl
- |
  prowler
- |
  proxemic
- |
  proxemics
- |
  proximal
- |
  proximally
- |
  proximate
- |
  proximately
- |
  proximation
- |
  proximity
- |
  proximo
- |
  proxy
- |
  Prozac
- |
  prude
- |
  Prudence
- |
  prudence
- |
  prudent
- |
  prudential
- |
  prudentially
- |
  prudently
- |
  prudery
- |
  prudish
- |
  prudishly
- |
  prudishness
- |
  prune
- |
  pruner
- |
  prurience
- |
  prurient
- |
  pruriently
- |
  Prussia
- |
  Prussian
- |
  pryer
- |
  pryingly
- |
  psalm
- |
  psalmist
- |
  psalmody
- |
  Psalms
- |
  Psalter
- |
  psalter
- |
  psaltery
- |
  psephologist
- |
  psephology
- |
  pseudo
- |
  pseudonym
- |
  pseudonymity
- |
  pseudonymous
- |
  pshaw
- |
  psittacosis
- |
  psoriasis
- |
  psych
- |
  Psyche
- |
  psyche
- |
  psyched
- |
  psychedelic
- |
  psychiatric
- |
  psychiatrist
- |
  psychiatry
- |
  psychic
- |
  psychical
- |
  psychically
- |
  psychics
- |
  psychism
- |
  psycho
- |
  psychoactive
- |
  psychobabble
- |
  psychodrama
- |
  psychogenic
- |
  psychologist
- |
  psychology
- |
  psychometry
- |
  psychomotor
- |
  psychopath
- |
  psychopathic
- |
  psychopathy
- |
  psychoses
- |
  psychosexual
- |
  psychosis
- |
  psychotic
- |
  psychotropic
- |
  ptarmigan
- |
  pterodactyl
- |
  pterosaur
- |
  Ptolemaic
- |
  Ptolemy
- |
  ptomaine
- |
  pubertal
- |
  puberty
- |
  pubes
- |
  pubescence
- |
  pubescent
- |
  pubic
- |
  pubis
- |
  public
- |
  publican
- |
  publication
- |
  publicise
- |
  publicist
- |
  publicity
- |
  publicize
- |
  publicly
- |
  publish
- |
  publishable
- |
  publisher
- |
  publishing
- |
  Puccini
- |
  pucker
- |
  puckered
- |
  puckish
- |
  puckishly
- |
  puckishness
- |
  pudding
- |
  puddinglike
- |
  puddle
- |
  puddling
- |
  pudenda
- |
  pudendum
- |
  pudginess
- |
  pudgy
- |
  Puebla
- |
  Pueblo
- |
  pueblo
- |
  puerile
- |
  puerilely
- |
  puerility
- |
  puerperal
- |
  puerperium
- |
  puffball
- |
  puffer
- |
  puffery
- |
  puffin
- |
  puffiness
- |
  puffy
- |
  pugilism
- |
  pugilist
- |
  pugilistic
- |
  pugnacious
- |
  pugnaciously
- |
  pugnacity
- |
  puissance
- |
  puissant
- |
  puissantly
- |
  pukka
- |
  Pulaski
- |
  pulchritude
- |
  puler
- |
  puling
- |
  Pulitzer
- |
  pullback
- |
  puller
- |
  pullet
- |
  pulley
- |
  Pullman
- |
  pullout
- |
  pullover
- |
  pullulate
- |
  pullulating
- |
  pullulation
- |
  pullup
- |
  pulmonary
- |
  pulmotor
- |
  pulpiness
- |
  pulpit
- |
  pulpwood
- |
  pulpy
- |
  pulsar
- |
  pulsate
- |
  pulsatile
- |
  pulsating
- |
  pulsation
- |
  pulsator
- |
  pulsatory
- |
  pulse
- |
  pulverize
- |
  pumice
- |
  pummel
- |
  pumper
- |
  pumpernickel
- |
  pumpkin
- |
  Punch
- |
  punch
- |
  puncheon
- |
  puncher
- |
  punchy
- |
  punctilio
- |
  punctilious
- |
  punctual
- |
  punctuality
- |
  punctually
- |
  punctuate
- |
  punctuation
- |
  puncture
- |
  pundit
- |
  punditry
- |
  pungency
- |
  pungent
- |
  pungently
- |
  Punic
- |
  punily
- |
  puniness
- |
  punish
- |
  punishable
- |
  punishing
- |
  punishment
- |
  punitive
- |
  punitively
- |
  punitiveness
- |
  Punjab
- |
  Punjabi
- |
  punkin
- |
  punning
- |
  punster
- |
  punter
- |
  punting
- |
  pupae
- |
  pupal
- |
  pupil
- |
  puppet
- |
  puppeteer
- |
  puppetry
- |
  Puppis
- |
  puppy
- |
  purblind
- |
  purblindness
- |
  purchasable
- |
  purchase
- |
  purchaser
- |
  purdah
- |
  purebred
- |
  puree
- |
  purely
- |
  pureness
- |
  purgation
- |
  purgative
- |
  purgatorial
- |
  purgatory
- |
  purge
- |
  purger
- |
  purging
- |
  purification
- |
  purificatory
- |
  purifier
- |
  purify
- |
  Purim
- |
  purine
- |
  purism
- |
  purist
- |
  puristic
- |
  Puritan
- |
  puritan
- |
  puritanical
- |
  Puritanism
- |
  puritanism
- |
  purity
- |
  purlieu
- |
  purlieus
- |
  purlieux
- |
  purloin
- |
  purloiner
- |
  purple
- |
  purplish
- |
  purport
- |
  purported
- |
  purportedly
- |
  purpose
- |
  purposeful
- |
  purposefully
- |
  purposeless
- |
  purposely
- |
  purposive
- |
  purposively
- |
  purse
- |
  purser
- |
  purslane
- |
  pursuance
- |
  pursuant
- |
  pursue
- |
  pursuer
- |
  pursuit
- |
  pursuivant
- |
  purulence
- |
  purulent
- |
  purvey
- |
  purveyance
- |
  purveyor
- |
  purview
- |
  Pusan
- |
  pushbutton
- |
  pushcart
- |
  pusher
- |
  pushily
- |
  pushiness
- |
  pushing
- |
  Pushkin
- |
  pushover
- |
  Pushtu
- |
  pushup
- |
  pushy
- |
  pussy
- |
  pussycat
- |
  pussyfoot
- |
  pustular
- |
  pustulate
- |
  pustule
- |
  putative
- |
  putatively
- |
  putdown
- |
  Putin
- |
  putout
- |
  putrefaction
- |
  putrefactive
- |
  putrefy
- |
  putrescence
- |
  putrescent
- |
  putrid
- |
  putridity
- |
  putridness
- |
  putsch
- |
  puttee
- |
  putter
- |
  putterer
- |
  putty
- |
  Putumayo
- |
  puzzle
- |
  puzzled
- |
  puzzlement
- |
  puzzler
- |
  puzzling
- |
  Pygmalion
- |
  pygmean
- |
  Pygmy
- |
  pygmy
- |
  pyjamas
- |
  pylon
- |
  pylori
- |
  pyloric
- |
  pylorus
- |
  Pyongyang
- |
  pyorrhea
- |
  pyorrheal
- |
  pyorrhoea
- |
  pyramid
- |
  pyramidal
- |
  pyramidally
- |
  pyramidical
- |
  Pyrenean
- |
  Pyrenees
- |
  pyrethrum
- |
  pyretic
- |
  Pyrex
- |
  pyrimidine
- |
  pyrite
- |
  pyrites
- |
  pyritic
- |
  pyrolysis
- |
  pyrolytic
- |
  pyromania
- |
  pyromaniac
- |
  pyromaniacal
- |
  pyromanic
- |
  pyrotechnic
- |
  pyrotechnics
- |
  pyrotechnist
- |
  Pyrrhic
- |
  pyrrhic
- |
  Pythagoras
- |
  Pythagorean
- |
  python
- |
  pythoness
- |
  Pyxis
- |
  Qabalah
- |
  Qaddafi
- |
  Qadhafi
- |
  Qatar
- |
  Qatari
- |
  qindarka
- |
  Qingdao
- |
  qintar
- |
  Qiqihar
- |
  qiviut
- |
  quack
- |
  quackery
- |
  quackish
- |
  quadrangle
- |
  quadrangular
- |
  quadrant
- |
  quadrantal
- |
  quadraphonic
- |
  quadratic
- |
  quadrennia
- |
  quadrennial
- |
  quadrennium
- |
  quadriceps
- |
  quadrille
- |
  quadrillion
- |
  quadriphonic
- |
  quadriplegia
- |
  quadriplegic
- |
  quadrivia
- |
  quadrivium
- |
  quadroon
- |
  quadruped
- |
  quadrupedal
- |
  quadruple
- |
  quadruplet
- |
  quaff
- |
  quaffer
- |
  quagmire
- |
  quahaug
- |
  quahog
- |
  quail
- |
  quaint
- |
  quaintly
- |
  quaintness
- |
  quake
- |
  Quaker
- |
  Quakerism
- |
  quaky
- |
  quale
- |
  qualia
- |
  qualified
- |
  qualifier
- |
  qualify
- |
  qualitative
- |
  quality
- |
  qualm
- |
  qualmish
- |
  quandary
- |
  quanta
- |
  quantifiable
- |
  quantifier
- |
  quantify
- |
  quantitative
- |
  quantities
- |
  quantity
- |
  quantize
- |
  quantum
- |
  quarantine
- |
  quark
- |
  quarrel
- |
  quarreler
- |
  quarreller
- |
  quarrelsome
- |
  quarrier
- |
  quarry
- |
  quarrying
- |
  quart
- |
  Quarter
- |
  quarter
- |
  quarterback
- |
  quarterdeck
- |
  quarterfinal
- |
  quarterly
- |
  quarters
- |
  quarterstaff
- |
  quartet
- |
  quartette
- |
  quartile
- |
  quarto
- |
  quartz
- |
  quartzite
- |
  quasar
- |
  quash
- |
  quasi
- |
  Quaternary
- |
  quaternary
- |
  quatrain
- |
  quatrefoil
- |
  quattrocento
- |
  quaver
- |
  quaveringly
- |
  quavery
- |
  Quayle
- |
  quean
- |
  queasily
- |
  queasiness
- |
  queasy
- |
  Quebec
- |
  Quebecer
- |
  Quebecker
- |
  Quebecois
- |
  Quechua
- |
  Quechuan
- |
  Queen
- |
  queen
- |
  queendom
- |
  queenlike
- |
  queenliness
- |
  queenly
- |
  Queens
- |
  queenship
- |
  Queensland
- |
  Queenslander
- |
  queer
- |
  queerly
- |
  queerness
- |
  quell
- |
  queller
- |
  Quemoy
- |
  quench
- |
  quenchable
- |
  quencher
- |
  quenchless
- |
  Quentin
- |
  Queretaro
- |
  querist
- |
  querulous
- |
  querulously
- |
  query
- |
  quesadilla
- |
  quest
- |
  quester
- |
  question
- |
  questionable
- |
  questionably
- |
  questioner
- |
  questioning
- |
  quetzal
- |
  Quetzalcoatl
- |
  queue
- |
  quibble
- |
  quibbler
- |
  quibbling
- |
  quiche
- |
  quick
- |
  quicken
- |
  quickie
- |
  quicklime
- |
  quickly
- |
  quickness
- |
  quicksand
- |
  quicksilver
- |
  quickstep
- |
  quiddity
- |
  quidnunc
- |
  quiescence
- |
  quiescent
- |
  quiescently
- |
  quiet
- |
  quietly
- |
  quietness
- |
  quietude
- |
  quietus
- |
  quill
- |
  Quilmes
- |
  quilt
- |
  quilted
- |
  quilter
- |
  quilting
- |
  quince
- |
  quinine
- |
  quinquennial
- |
  quinsy
- |
  quint
- |
  quintal
- |
  quintessence
- |
  quintet
- |
  quintette
- |
  quintile
- |
  Quintilian
- |
  quintillion
- |
  Quintin
- |
  quintuple
- |
  quintuplet
- |
  quipster
- |
  quire
- |
  quirk
- |
  quirkiness
- |
  quirkish
- |
  quirky
- |
  quirt
- |
  Quisling
- |
  quisling
- |
  quitclaim
- |
  quite
- |
  Quito
- |
  quits
- |
  quittance
- |
  quitter
- |
  quiver
- |
  quiveringly
- |
  quivery
- |
  quixotic
- |
  quixotically
- |
  quixotism
- |
  quixotry
- |
  quizzer
- |
  quizzical
- |
  quizzicality
- |
  quizzically
- |
  quodlibet
- |
  quoin
- |
  quoit
- |
  quoits
- |
  quondam
- |
  quorum
- |
  quota
- |
  quotability
- |
  quotable
- |
  quotation
- |
  quote
- |
  quoter
- |
  quoth
- |
  quotidian
- |
  quotient
- |
  qwerty
- |
  Rabat
- |
  rabbet
- |
  rabbi
- |
  rabbinate
- |
  rabbinic
- |
  rabbinical
- |
  rabbinically
- |
  rabbit
- |
  rabble
- |
  Rabelais
- |
  Rabelaisian
- |
  Rabia
- |
  rabid
- |
  rabidity
- |
  rabidly
- |
  rabidness
- |
  rabies
- |
  Rabin
- |
  raccoon
- |
  racecourse
- |
  racehorse
- |
  raceme
- |
  racemose
- |
  racer
- |
  races
- |
  racetrack
- |
  raceway
- |
  Rachel
- |
  rachitic
- |
  rachitis
- |
  Rachmaninoff
- |
  racial
- |
  racialism
- |
  racialist
- |
  racialistic
- |
  racialize
- |
  racially
- |
  racily
- |
  Racine
- |
  raciness
- |
  racing
- |
  racism
- |
  racist
- |
  racket
- |
  racketball
- |
  racketeer
- |
  racketeering
- |
  raconteur
- |
  raconteuse
- |
  racquet
- |
  racquetball
- |
  radar
- |
  radarscope
- |
  radial
- |
  radially
- |
  radian
- |
  radiance
- |
  radiancy
- |
  radiant
- |
  radiantly
- |
  radiate
- |
  radiation
- |
  radiational
- |
  radiative
- |
  radiator
- |
  radical
- |
  radicalism
- |
  radicalize
- |
  radically
- |
  radicalness
- |
  radicchio
- |
  radii
- |
  radio
- |
  radioactive
- |
  radiocarbon
- |
  radiogram
- |
  radiograph
- |
  radiographer
- |
  radiographic
- |
  radiography
- |
  radioisotope
- |
  radiologic
- |
  radiological
- |
  radiologist
- |
  radiology
- |
  radioman
- |
  radiometer
- |
  radiometric
- |
  radiometry
- |
  radiopacity
- |
  radiopaque
- |
  radiophone
- |
  radiophonic
- |
  radioscopic
- |
  radioscopy
- |
  radiosonde
- |
  radiotherapy
- |
  radish
- |
  radium
- |
  radius
- |
  radon
- |
  Rafael
- |
  raffia
- |
  raffish
- |
  raffishly
- |
  raffishness
- |
  raffle
- |
  rafter
- |
  rafting
- |
  ragamuffin
- |
  ragbag
- |
  ragged
- |
  raggedly
- |
  raggedness
- |
  raggedy
- |
  raging
- |
  ragingly
- |
  raglan
- |
  ragout
- |
  ragpicker
- |
  ragtag
- |
  ragtime
- |
  ragtop
- |
  ragweed
- |
  raider
- |
  railer
- |
  railing
- |
  raillery
- |
  railroad
- |
  railroader
- |
  railroading
- |
  railway
- |
  raiment
- |
  rainbow
- |
  raincoat
- |
  raindrop
- |
  rainfall
- |
  rainforest
- |
  Rainier
- |
  raininess
- |
  rainmaker
- |
  rainmaking
- |
  rainproof
- |
  rains
- |
  rainstorm
- |
  rainwater
- |
  rainy
- |
  raise
- |
  raiser
- |
  raisin
- |
  Rajab
- |
  rajah
- |
  Rajasthan
- |
  Rajkot
- |
  Rajputana
- |
  Rajshahi
- |
  raker
- |
  rakish
- |
  rakishly
- |
  rakishness
- |
  Ralegh
- |
  Raleigh
- |
  rales
- |
  rallier
- |
  rally
- |
  Ralph
- |
  Ramadan
- |
  ramble
- |
  rambler
- |
  rambling
- |
  rambunctious
- |
  ramekin
- |
  ramen
- |
  ramequin
- |
  Rameses
- |
  Ramesses
- |
  ramie
- |
  ramification
- |
  ramify
- |
  ramjet
- |
  Ramon
- |
  Ramona
- |
  rampage
- |
  rampageous
- |
  rampager
- |
  rampancy
- |
  rampant
- |
  rampantly
- |
  rampart
- |
  ramrod
- |
  Ramsay
- |
  Ramses
- |
  ramshackle
- |
  ranch
- |
  rancher
- |
  rancheria
- |
  ranchero
- |
  Ranchi
- |
  ranching
- |
  rancho
- |
  rancid
- |
  rancidity
- |
  rancidness
- |
  rancor
- |
  rancorous
- |
  rancorously
- |
  rancour
- |
  Randal
- |
  Randall
- |
  randiness
- |
  Randolph
- |
  random
- |
  randomize
- |
  randomly
- |
  randomness
- |
  Randwick
- |
  Randy
- |
  randy
- |
  ranee
- |
  range
- |
  Ranger
- |
  ranger
- |
  ranginess
- |
  Rangoon
- |
  rangy
- |
  Rankin
- |
  ranking
- |
  rankle
- |
  rankly
- |
  rankness
- |
  ranks
- |
  ransack
- |
  ransacking
- |
  ransom
- |
  ransomer
- |
  ranter
- |
  ranting
- |
  rantingly
- |
  rapacious
- |
  rapaciously
- |
  rapacity
- |
  raper
- |
  rapeseed
- |
  Raphael
- |
  rapid
- |
  rapidity
- |
  rapidly
- |
  rapidness
- |
  rapids
- |
  rapier
- |
  rapine
- |
  rapist
- |
  rappel
- |
  rappen
- |
  rapper
- |
  rapport
- |
  rapporteur
- |
  rapscallion
- |
  raptly
- |
  raptness
- |
  raptor
- |
  raptorial
- |
  raptorially
- |
  Rapture
- |
  rapture
- |
  raptures
- |
  rapturous
- |
  rapturously
- |
  rarebit
- |
  rarefaction
- |
  rarefiable
- |
  rarefied
- |
  rarefy
- |
  rarely
- |
  rareness
- |
  rarified
- |
  rarify
- |
  raring
- |
  rarity
- |
  Rasalgethi
- |
  Rasalhague
- |
  rascal
- |
  rascality
- |
  rascally
- |
  rasher
- |
  rashly
- |
  rashness
- |
  Rasht
- |
  raspberry
- |
  raspiness
- |
  Rasputin
- |
  raspy
- |
  Rastafarian
- |
  raster
- |
  ratatouille
- |
  ratchet
- |
  rater
- |
  Rathaus
- |
  Rathauser
- |
  rathe
- |
  rather
- |
  rathskeller
- |
  ratifiable
- |
  ratification
- |
  ratifier
- |
  ratify
- |
  rating
- |
  ratings
- |
  ratio
- |
  ratiocinate
- |
  ratiocinator
- |
  ration
- |
  rational
- |
  rationale
- |
  rationalise
- |
  rationalism
- |
  rationalist
- |
  rationality
- |
  rationalize
- |
  rationalizer
- |
  rationally
- |
  rationalness
- |
  rationing
- |
  rations
- |
  ratlike
- |
  ratlin
- |
  ratline
- |
  rattan
- |
  ratter
- |
  rattiness
- |
  rattle
- |
  rattlebrain
- |
  rattled
- |
  rattler
- |
  rattlesnake
- |
  rattletrap
- |
  rattling
- |
  rattly
- |
  rattrap
- |
  ratty
- |
  raucous
- |
  raucously
- |
  raucousness
- |
  raunchily
- |
  raunchiness
- |
  raunchy
- |
  ravage
- |
  ravager
- |
  ravages
- |
  Ravel
- |
  ravel
- |
  raveler
- |
  raveling
- |
  ravelling
- |
  raven
- |
  ravening
- |
  Ravenna
- |
  ravenous
- |
  ravenously
- |
  ravenousness
- |
  ravine
- |
  raving
- |
  ravingly
- |
  ravings
- |
  ravioli
- |
  ravish
- |
  ravisher
- |
  ravishing
- |
  ravishingly
- |
  ravishment
- |
  Rawalpindi
- |
  rawboned
- |
  rawhide
- |
  Rawlings
- |
  rawness
- |
  Raymond
- |
  rayon
- |
  razor
- |
  razorback
- |
  razzmatazz
- |
  reabsorb
- |
  reabsorption
- |
  reach
- |
  reachable
- |
  reacher
- |
  reaches
- |
  reacquaint
- |
  reacquire
- |
  react
- |
  reactance
- |
  reactant
- |
  reaction
- |
  reactionary
- |
  reactions
- |
  reactivate
- |
  reactivation
- |
  reactive
- |
  reactivity
- |
  reactor
- |
  readability
- |
  readable
- |
  readableness
- |
  readably
- |
  readapt
- |
  readdress
- |
  reader
- |
  readership
- |
  readily
- |
  readiness
- |
  Reading
- |
  reading
- |
  readjourn
- |
  readjust
- |
  readjustment
- |
  readmission
- |
  readmit
- |
  readmittance
- |
  readopt
- |
  readoption
- |
  readout
- |
  ready
- |
  reaffirm
- |
  Reagan
- |
  reagent
- |
  realign
- |
  realignment
- |
  realise
- |
  realism
- |
  realist
- |
  realistic
- |
  reality
- |
  realizable
- |
  realization
- |
  realize
- |
  reallocate
- |
  reallocation
- |
  really
- |
  realm
- |
  realness
- |
  realpolitik
- |
  Realtor
- |
  realtor
- |
  realty
- |
  reamer
- |
  reams
- |
  reanalysis
- |
  reanalyze
- |
  reanimate
- |
  reanimation
- |
  reannex
- |
  reannexation
- |
  reaper
- |
  reappear
- |
  reappearance
- |
  reapply
- |
  reappoint
- |
  reapportion
- |
  reappraisal
- |
  reappraise
- |
  rearguard
- |
  rearm
- |
  rearmament
- |
  rearmost
- |
  rearouse
- |
  rearrange
- |
  rearrest
- |
  rearward
- |
  rearwards
- |
  reascend
- |
  reason
- |
  reasonable
- |
  reasonably
- |
  reasoned
- |
  reasoner
- |
  reasoning
- |
  reassemble
- |
  reassembly
- |
  reassert
- |
  reassertion
- |
  reassess
- |
  reassessment
- |
  reassign
- |
  reassignment
- |
  reassume
- |
  reassurance
- |
  reassure
- |
  reassured
- |
  reassuring
- |
  reassuringly
- |
  reattach
- |
  reattachment
- |
  reattain
- |
  reattainment
- |
  reattempt
- |
  reauthorize
- |
  reave
- |
  reaver
- |
  reawake
- |
  reawaken
- |
  reawoke
- |
  rebaptism
- |
  rebaptize
- |
  rebarbative
- |
  rebatable
- |
  rebate
- |
  rebater
- |
  Rebecca
- |
  Rebekah
- |
  rebel
- |
  rebellion
- |
  rebellious
- |
  rebelliously
- |
  rebid
- |
  rebind
- |
  rebirth
- |
  reboil
- |
  reboot
- |
  reborn
- |
  rebound
- |
  rebroadcast
- |
  rebuff
- |
  rebuild
- |
  rebuilt
- |
  rebuke
- |
  rebukingly
- |
  reburial
- |
  rebury
- |
  rebus
- |
  rebut
- |
  rebuttable
- |
  rebuttal
- |
  rebutter
- |
  recalcitrant
- |
  recalculate
- |
  recall
- |
  recant
- |
  recantation
- |
  recanter
- |
  recap
- |
  recapitalize
- |
  recapitulate
- |
  recapture
- |
  recast
- |
  recede
- |
  receding
- |
  receipt
- |
  receipts
- |
  receivable
- |
  receivables
- |
  receive
- |
  received
- |
  receiver
- |
  receivership
- |
  recency
- |
  recension
- |
  recent
- |
  recently
- |
  recentness
- |
  receptacle
- |
  reception
- |
  receptionist
- |
  receptive
- |
  receptively
- |
  receptivity
- |
  receptor
- |
  recess
- |
  recesses
- |
  recession
- |
  recessional
- |
  recessionary
- |
  recessive
- |
  recessively
- |
  recessivity
- |
  rechannel
- |
  recharge
- |
  rechargeable
- |
  recharter
- |
  recheck
- |
  recherche
- |
  rechristen
- |
  recidivism
- |
  recidivist
- |
  recidivistic
- |
  recidivous
- |
  Recife
- |
  recipe
- |
  recipient
- |
  reciprocal
- |
  reciprocally
- |
  reciprocate
- |
  reciprocator
- |
  reciprocity
- |
  recirculate
- |
  recital
- |
  recitalist
- |
  recitation
- |
  recitative
- |
  recite
- |
  reciter
- |
  reckless
- |
  recklessly
- |
  recklessness
- |
  reckon
- |
  reckoning
- |
  reclaim
- |
  reclaimable
- |
  reclaimant
- |
  reclaimer
- |
  reclamation
- |
  reclassify
- |
  recline
- |
  recliner
- |
  reclothe
- |
  recluse
- |
  reclusion
- |
  reclusive
- |
  recognisable
- |
  recognise
- |
  recognition
- |
  recognizable
- |
  recognizably
- |
  recognizance
- |
  recognizant
- |
  recognize
- |
  recoil
- |
  recoilless
- |
  recoin
- |
  recollect
- |
  recollection
- |
  recolonize
- |
  recolor
- |
  recomb
- |
  recombine
- |
  recommence
- |
  recommend
- |
  recommended
- |
  recommission
- |
  recommit
- |
  recommitment
- |
  recompense
- |
  recompile
- |
  recompose
- |
  recompute
- |
  reconceive
- |
  reconception
- |
  reconcilable
- |
  reconcile
- |
  reconciled
- |
  reconciler
- |
  recondense
- |
  recondite
- |
  recondition
- |
  reconduct
- |
  reconfirm
- |
  reconnect
- |
  reconnection
- |
  reconnoiter
- |
  reconnoitre
- |
  reconquer
- |
  reconquest
- |
  reconsecrate
- |
  reconsider
- |
  reconsign
- |
  reconstitute
- |
  reconstruct
- |
  recontact
- |
  recontract
- |
  reconvene
- |
  reconversion
- |
  reconvert
- |
  reconvey
- |
  recook
- |
  recopy
- |
  record
- |
  recorder
- |
  recording
- |
  recordist
- |
  recount
- |
  recoup
- |
  recoupable
- |
  recoupment
- |
  recourse
- |
  recover
- |
  recoverable
- |
  recovery
- |
  recreance
- |
  recreancy
- |
  recreant
- |
  recreantly
- |
  recreate
- |
  recreation
- |
  recreational
- |
  recreative
- |
  recriminate
- |
  recross
- |
  recrudesce
- |
  recrudescent
- |
  recruit
- |
  recruiter
- |
  recruiting
- |
  recruitment
- |
  recta
- |
  rectal
- |
  rectally
- |
  rectangle
- |
  rectangular
- |
  rectifiable
- |
  rectified
- |
  rectifier
- |
  rectify
- |
  rectilineal
- |
  rectilinear
- |
  rectitude
- |
  recto
- |
  rector
- |
  rectorate
- |
  rectorial
- |
  rectorship
- |
  rectory
- |
  rectum
- |
  recumbency
- |
  recumbent
- |
  recumbently
- |
  recuperable
- |
  recuperate
- |
  recuperation
- |
  recuperative
- |
  recur
- |
  recurrence
- |
  recurrent
- |
  recurrently
- |
  recursive
- |
  recursively
- |
  recurvature
- |
  recurve
- |
  recusal
- |
  recusance
- |
  recusancy
- |
  recusant
- |
  recuse
- |
  recut
- |
  recyclable
- |
  recycle
- |
  recycled
- |
  recycler
- |
  recycling
- |
  redact
- |
  redaction
- |
  redactor
- |
  redbreast
- |
  Redbridge
- |
  redcap
- |
  redcoat
- |
  redden
- |
  reddish
- |
  reddishness
- |
  redecorate
- |
  redecoration
- |
  rededicate
- |
  rededication
- |
  redeem
- |
  redeemable
- |
  redeemer
- |
  redeeming
- |
  redefine
- |
  redefinition
- |
  redeliver
- |
  redemption
- |
  redemptional
- |
  redemptive
- |
  redemptory
- |
  redeploy
- |
  redeployment
- |
  redeposit
- |
  redesign
- |
  redetermine
- |
  redevelop
- |
  Redgrave
- |
  redhead
- |
  redheaded
- |
  redial
- |
  redid
- |
  redigest
- |
  redintegrate
- |
  redirect
- |
  redirection
- |
  rediscount
- |
  rediscover
- |
  rediscovery
- |
  redissolve
- |
  redistill
- |
  redistribute
- |
  redistrict
- |
  redivide
- |
  redivivus
- |
  redline
- |
  redlining
- |
  redly
- |
  redneck
- |
  redness
- |
  redolence
- |
  redolent
- |
  redolently
- |
  redone
- |
  redouble
- |
  redoubt
- |
  redoubtable
- |
  redoubtably
- |
  redound
- |
  redraft
- |
  redraw
- |
  redrawn
- |
  redress
- |
  redressable
- |
  redressal
- |
  redresser
- |
  redrew
- |
  redshift
- |
  reduce
- |
  reducer
- |
  reducibility
- |
  reducible
- |
  reduction
- |
  reductive
- |
  redundancy
- |
  redundant
- |
  redundantly
- |
  reduplicate
- |
  redux
- |
  redwood
- |
  redye
- |
  reecho
- |
  reediness
- |
  reedit
- |
  reeducate
- |
  reeducation
- |
  reedy
- |
  reefer
- |
  reeker
- |
  reeky
- |
  reelable
- |
  reelect
- |
  reelection
- |
  reeler
- |
  reembark
- |
  reembody
- |
  reemerge
- |
  reemergence
- |
  reemphasis
- |
  reemphasize
- |
  reemploy
- |
  reemployment
- |
  reenact
- |
  reenactment
- |
  reenergize
- |
  reengage
- |
  reenlist
- |
  reenlistment
- |
  reenter
- |
  reentrance
- |
  reentry
- |
  reequip
- |
  reestablish
- |
  reevaluate
- |
  reevaluation
- |
  reeve
- |
  reexamine
- |
  reexchange
- |
  reexhibit
- |
  reexperience
- |
  reexplain
- |
  reexport
- |
  reface
- |
  refashion
- |
  refasten
- |
  refection
- |
  refectory
- |
  refer
- |
  referable
- |
  referee
- |
  reference
- |
  referenda
- |
  referendum
- |
  referent
- |
  referential
- |
  referral
- |
  referrer
- |
  refight
- |
  refile
- |
  refill
- |
  refillable
- |
  refilm
- |
  refilter
- |
  refinance
- |
  refine
- |
  refined
- |
  refinement
- |
  refiner
- |
  refinery
- |
  refining
- |
  refinish
- |
  refinisher
- |
  refire
- |
  refit
- |
  refix
- |
  reflect
- |
  reflection
- |
  reflective
- |
  reflectively
- |
  reflectivity
- |
  reflector
- |
  reflex
- |
  reflexion
- |
  reflexive
- |
  reflexively
- |
  reflexivity
- |
  reflexly
- |
  reflexology
- |
  refloat
- |
  reflow
- |
  reflower
- |
  reflux
- |
  refocus
- |
  refold
- |
  reforest
- |
  reforge
- |
  reform
- |
  reformable
- |
  reformat
- |
  Reformation
- |
  reformation
- |
  reformative
- |
  reformatory
- |
  reformed
- |
  reformer
- |
  reformist
- |
  reformulate
- |
  refortify
- |
  refound
- |
  refract
- |
  refraction
- |
  refractional
- |
  refractive
- |
  refractively
- |
  refractivity
- |
  refractor
- |
  refractorily
- |
  refractory
- |
  refrain
- |
  refrainment
- |
  refreeze
- |
  refresh
- |
  refreshed
- |
  refresher
- |
  refreshing
- |
  refreshingly
- |
  refreshment
- |
  refreshments
- |
  refrigerant
- |
  refrigerate
- |
  refrigerator
- |
  refroze
- |
  refrozen
- |
  refry
- |
  refuel
- |
  refueling
- |
  refuelling
- |
  refuge
- |
  refugee
- |
  refulgence
- |
  refulgent
- |
  refulgently
- |
  refund
- |
  refundable
- |
  refurbish
- |
  refurnish
- |
  refusal
- |
  refuse
- |
  refutable
- |
  refutably
- |
  refutal
- |
  refutation
- |
  refute
- |
  refuter
- |
  regain
- |
  regal
- |
  regale
- |
  regalement
- |
  regalia
- |
  regality
- |
  regally
- |
  regard
- |
  regardful
- |
  regarding
- |
  regardless
- |
  regardlessly
- |
  regards
- |
  regather
- |
  regatta
- |
  regear
- |
  Regency
- |
  regency
- |
  regeneracy
- |
  regenerate
- |
  regeneration
- |
  regenerative
- |
  regenerator
- |
  regent
- |
  regerminate
- |
  reggae
- |
  Reggie
- |
  regicidal
- |
  regicide
- |
  regild
- |
  regime
- |
  regimen
- |
  regiment
- |
  regimental
- |
  regimentals
- |
  regimented
- |
  Regina
- |
  Reginald
- |
  region
- |
  regional
- |
  regionalism
- |
  regionally
- |
  Regis
- |
  regisseur
- |
  register
- |
  registered
- |
  registrable
- |
  registrant
- |
  registrar
- |
  registration
- |
  registry
- |
  regive
- |
  reglaze
- |
  regnant
- |
  regolith
- |
  regrade
- |
  regress
- |
  regression
- |
  regressive
- |
  regressively
- |
  regressor
- |
  regret
- |
  regretful
- |
  regretfully
- |
  regrets
- |
  regrettable
- |
  regrettably
- |
  regretter
- |
  regrew
- |
  regrind
- |
  regroup
- |
  regrow
- |
  regrown
- |
  regrowth
- |
  regular
- |
  regularity
- |
  regularize
- |
  regularly
- |
  regulate
- |
  regulated
- |
  regulation
- |
  regulative
- |
  regulator
- |
  regulatory
- |
  Regulus
- |
  regurgitate
- |
  rehab
- |
  rehabilitate
- |
  rehandle
- |
  rehang
- |
  rehash
- |
  rehear
- |
  rehearing
- |
  rehearsal
- |
  rehearse
- |
  rehearser
- |
  reheat
- |
  rehire
- |
  Rehnquist
- |
  rehouse
- |
  rehung
- |
  Reich
- |
  reification
- |
  reificatory
- |
  reify
- |
  reign
- |
  reigning
- |
  reignite
- |
  reimbursable
- |
  reimburse
- |
  reimport
- |
  reimpose
- |
  reimposition
- |
  reimpress
- |
  reimprison
- |
  Reims
- |
  reincarnate
- |
  reincur
- |
  reindeer
- |
  reinduce
- |
  reinfect
- |
  reinfection
- |
  reinflame
- |
  reinforce
- |
  reinforced
- |
  reinforcer
- |
  reinfuse
- |
  reinfusion
- |
  reinoculate
- |
  reins
- |
  reinscribe
- |
  reinsert
- |
  reinsertion
- |
  reinspect
- |
  reinstate
- |
  reinstruct
- |
  reinsure
- |
  reintegrate
- |
  reinter
- |
  reinterpret
- |
  reintroduce
- |
  reinvent
- |
  reinvention
- |
  reinvest
- |
  reinvestment
- |
  reinvigorate
- |
  reissue
- |
  reiterate
- |
  reiteration
- |
  reiterative
- |
  reject
- |
  rejecter
- |
  rejection
- |
  rejoice
- |
  rejoicer
- |
  rejoicing
- |
  rejoin
- |
  rejoinder
- |
  rejudge
- |
  rejuvenate
- |
  rejuvenated
- |
  rejuvenating
- |
  rejuvenation
- |
  rejuvenator
- |
  rekindle
- |
  reknit
- |
  relabel
- |
  relaid
- |
  relapse
- |
  relapser
- |
  relatable
- |
  relate
- |
  related
- |
  relatedness
- |
  relater
- |
  relation
- |
  relational
- |
  relations
- |
  relationship
- |
  relative
- |
  relatively
- |
  relativeness
- |
  relativism
- |
  relativist
- |
  relativistic
- |
  relativity
- |
  relator
- |
  relaunch
- |
  relax
- |
  relaxant
- |
  relaxation
- |
  relaxed
- |
  relaxer
- |
  relaxing
- |
  relay
- |
  relearn
- |
  releasable
- |
  release
- |
  releaser
- |
  relegate
- |
  relegation
- |
  relent
- |
  relentless
- |
  relentlessly
- |
  relevance
- |
  relevancy
- |
  relevant
- |
  relevantly
- |
  reliability
- |
  reliable
- |
  reliableness
- |
  reliably
- |
  reliance
- |
  reliant
- |
  reliantly
- |
  relic
- |
  relics
- |
  relict
- |
  relief
- |
  relieve
- |
  relieved
- |
  reliever
- |
  relight
- |
  religion
- |
  religionist
- |
  religiose
- |
  religiosity
- |
  religious
- |
  religiously
- |
  reline
- |
  relinquish
- |
  relinquisher
- |
  reliquary
- |
  reliquiae
- |
  relish
- |
  relishable
- |
  relivable
- |
  relive
- |
  reload
- |
  relocate
- |
  relocation
- |
  reluctance
- |
  reluctant
- |
  reluctantly
- |
  remade
- |
  remain
- |
  remainder
- |
  remaining
- |
  remains
- |
  remake
- |
  remand
- |
  remandment
- |
  remanence
- |
  remanent
- |
  remap
- |
  remark
- |
  remarkable
- |
  remarkably
- |
  Remarque
- |
  remarriage
- |
  remarry
- |
  rematch
- |
  Rembrandt
- |
  remeasure
- |
  remediable
- |
  remedial
- |
  remedially
- |
  remediless
- |
  remedy
- |
  remelt
- |
  remember
- |
  rememberable
- |
  remembrance
- |
  remigrate
- |
  remigration
- |
  remilitarize
- |
  remind
- |
  reminder
- |
  Remington
- |
  reminisce
- |
  reminiscence
- |
  reminiscent
- |
  remiss
- |
  remissible
- |
  remissibly
- |
  remission
- |
  remissly
- |
  remissness
- |
  remit
- |
  remittable
- |
  remittal
- |
  remittance
- |
  remittent
- |
  remitter
- |
  remix
- |
  remnant
- |
  remodel
- |
  remodeler
- |
  remodify
- |
  remold
- |
  remonetize
- |
  remonstrance
- |
  remonstrant
- |
  remonstrate
- |
  remonstrator
- |
  remora
- |
  remorse
- |
  remorseful
- |
  remorsefully
- |
  remorseless
- |
  remote
- |
  remotely
- |
  remoteness
- |
  remount
- |
  removable
- |
  removably
- |
  removal
- |
  remove
- |
  removed
- |
  remover
- |
  remunerate
- |
  remuneration
- |
  remunerative
- |
  remunerator
- |
  Remus
- |
  Renaissance
- |
  renaissance
- |
  renal
- |
  rename
- |
  Renascence
- |
  renascence
- |
  renascent
- |
  Renault
- |
  render
- |
  renderer
- |
  rendering
- |
  rendezvous
- |
  rendition
- |
  Renee
- |
  renegade
- |
  renege
- |
  reneger
- |
  renegotiate
- |
  renew
- |
  renewable
- |
  renewal
- |
  renewed
- |
  renewer
- |
  Rennes
- |
  rennet
- |
  rennin
- |
  Renoir
- |
  renominate
- |
  renomination
- |
  renotify
- |
  renounce
- |
  renounceable
- |
  renouncement
- |
  renouncer
- |
  renovate
- |
  renovation
- |
  renovator
- |
  renown
- |
  renowned
- |
  rentable
- |
  rental
- |
  renter
- |
  rentier
- |
  renumber
- |
  renunciant
- |
  renunciation
- |
  renunciative
- |
  renunciatory
- |
  reoccupation
- |
  reoccupy
- |
  reoccur
- |
  reoccurrence
- |
  reopen
- |
  reorder
- |
  reorganize
- |
  reorient
- |
  reorientate
- |
  repack
- |
  repackage
- |
  repaid
- |
  repaint
- |
  repair
- |
  repairable
- |
  repairer
- |
  repairman
- |
  repairwoman
- |
  reparable
- |
  reparably
- |
  reparation
- |
  reparations
- |
  reparative
- |
  reparatory
- |
  repartee
- |
  repass
- |
  repast
- |
  repatriate
- |
  repatriation
- |
  repave
- |
  repay
- |
  repayable
- |
  repayment
- |
  repeal
- |
  repealable
- |
  repealer
- |
  repeat
- |
  repeatable
- |
  repeated
- |
  repeatedly
- |
  repeater
- |
  repechage
- |
  repel
- |
  repellant
- |
  repelled
- |
  repellence
- |
  repellency
- |
  repellent
- |
  repellently
- |
  repent
- |
  repentance
- |
  repentant
- |
  repentantly
- |
  repenter
- |
  repeople
- |
  repercussion
- |
  repercussive
- |
  repertoire
- |
  repertorial
- |
  repertory
- |
  repetend
- |
  repetition
- |
  repetitious
- |
  repetitive
- |
  repetitively
- |
  rephotograph
- |
  rephrase
- |
  repine
- |
  repiner
- |
  replace
- |
  replaceable
- |
  replacement
- |
  replacer
- |
  replant
- |
  replay
- |
  replenish
- |
  replenisher
- |
  replete
- |
  repleteness
- |
  repletion
- |
  replevin
- |
  replica
- |
  replicable
- |
  replicate
- |
  replication
- |
  replicative
- |
  replier
- |
  reply
- |
  repopulate
- |
  report
- |
  reportable
- |
  reportage
- |
  reportedly
- |
  reporter
- |
  reporting
- |
  reportorial
- |
  repose
- |
  reposeful
- |
  reposefully
- |
  repository
- |
  repossess
- |
  repossession
- |
  repousse
- |
  reprehend
- |
  reprehension
- |
  represent
- |
  repress
- |
  repressed
- |
  represser
- |
  repressible
- |
  repression
- |
  repressive
- |
  repressively
- |
  repressor
- |
  reprice
- |
  reprieve
- |
  reprimand
- |
  reprint
- |
  reprinter
- |
  reprisal
- |
  reprise
- |
  reproach
- |
  reproachable
- |
  reproacher
- |
  reproachful
- |
  reprobate
- |
  reprobation
- |
  reprocess
- |
  reproduce
- |
  reproducer
- |
  reproducible
- |
  reproduction
- |
  reproductive
- |
  reprogram
- |
  reproof
- |
  reprovable
- |
  reproval
- |
  reprove
- |
  reprover
- |
  reprovingly
- |
  reptile
- |
  reptilian
- |
  republic
- |
  Republican
- |
  republican
- |
  republish
- |
  repudiate
- |
  repudiation
- |
  repudiator
- |
  repugnance
- |
  repugnant
- |
  repugnantly
- |
  repulse
- |
  repulsion
- |
  repulsive
- |
  repulsively
- |
  repurchase
- |
  reputability
- |
  reputable
- |
  reputably
- |
  reputation
- |
  repute
- |
  reputed
- |
  reputedly
- |
  request
- |
  requester
- |
  Requiem
- |
  requiem
- |
  require
- |
  required
- |
  requirement
- |
  requisite
- |
  requisitely
- |
  requisition
- |
  requitable
- |
  requital
- |
  requite
- |
  requiter
- |
  reradiate
- |
  reran
- |
  reread
- |
  rereading
- |
  rerecord
- |
  reredos
- |
  rerelease
- |
  reroute
- |
  rerun
- |
  resalable
- |
  resale
- |
  reschedule
- |
  rescheduling
- |
  rescind
- |
  rescindable
- |
  rescission
- |
  rescore
- |
  rescreen
- |
  rescript
- |
  rescue
- |
  rescuer
- |
  reseal
- |
  resealable
- |
  research
- |
  researcher
- |
  reseau
- |
  reseaux
- |
  resect
- |
  resected
- |
  resection
- |
  resectional
- |
  reseed
- |
  resegregate
- |
  resell
- |
  resemblance
- |
  resemble
- |
  resent
- |
  resentful
- |
  resentfully
- |
  resentment
- |
  reserpine
- |
  reservable
- |
  reservation
- |
  reserve
- |
  reserved
- |
  reservedly
- |
  reservedness
- |
  reserves
- |
  reservist
- |
  reservoir
- |
  reset
- |
  resettle
- |
  resettlement
- |
  resew
- |
  reshape
- |
  reshaping
- |
  resharpen
- |
  reship
- |
  reshipment
- |
  reshow
- |
  reshuffle
- |
  reside
- |
  residence
- |
  residency
- |
  resident
- |
  residential
- |
  residentship
- |
  resider
- |
  residua
- |
  residual
- |
  residually
- |
  residuals
- |
  residuary
- |
  residue
- |
  residuum
- |
  resign
- |
  resignation
- |
  resigned
- |
  resignedly
- |
  resilience
- |
  resiliency
- |
  resilient
- |
  resiliently
- |
  resin
- |
  resined
- |
  resinous
- |
  resist
- |
  Resistance
- |
  resistance
- |
  resistant
- |
  resister
- |
  resistible
- |
  resistless
- |
  resistor
- |
  resold
- |
  resole
- |
  resolute
- |
  resolutely
- |
  resoluteness
- |
  resolution
- |
  resolvable
- |
  resolve
- |
  resolved
- |
  resolver
- |
  resonance
- |
  resonant
- |
  resonantly
- |
  resonate
- |
  resonator
- |
  resorption
- |
  resort
- |
  resound
- |
  resounding
- |
  resoundingly
- |
  resource
- |
  resourceful
- |
  resources
- |
  resow
- |
  respect
- |
  respectable
- |
  respectably
- |
  respected
- |
  respecter
- |
  respectful
- |
  respectfully
- |
  respecting
- |
  respective
- |
  respectively
- |
  respects
- |
  respell
- |
  respiration
- |
  respirator
- |
  respiratory
- |
  respire
- |
  respite
- |
  resplendence
- |
  resplendency
- |
  resplendent
- |
  respond
- |
  respondent
- |
  responder
- |
  response
- |
  responsible
- |
  responsibly
- |
  responsive
- |
  responsively
- |
  respray
- |
  ressentiment
- |
  restack
- |
  restaff
- |
  restage
- |
  restart
- |
  restate
- |
  restatement
- |
  restaurant
- |
  restaurateur
- |
  rester
- |
  restful
- |
  restfully
- |
  restfulness
- |
  restitch
- |
  restitution
- |
  restitutive
- |
  restive
- |
  restively
- |
  restiveness
- |
  restless
- |
  restlessly
- |
  restlessness
- |
  restock
- |
  restorable
- |
  Restoration
- |
  restoration
- |
  restorative
- |
  restore
- |
  restorer
- |
  restraighten
- |
  restrain
- |
  restrainable
- |
  restrained
- |
  restrainedly
- |
  restrainer
- |
  restraining
- |
  restraint
- |
  restraints
- |
  restrengthen
- |
  restrict
- |
  restricted
- |
  restriction
- |
  restrictive
- |
  restrike
- |
  restring
- |
  restroom
- |
  restructure
- |
  restrung
- |
  restudy
- |
  restuff
- |
  restyle
- |
  resubmission
- |
  resubmit
- |
  resubscribe
- |
  result
- |
  resultant
- |
  results
- |
  resumable
- |
  resume
- |
  resummon
- |
  resumption
- |
  resumptive
- |
  resupply
- |
  resurface
- |
  resurgence
- |
  resurgent
- |
  resurrect
- |
  Resurrection
- |
  resurrection
- |
  resurvey
- |
  resuscitate
- |
  resuscitator
- |
  resynthesis
- |
  resynthesize
- |
  retable
- |
  retablo
- |
  retail
- |
  retailer
- |
  retailing
- |
  retain
- |
  retainable
- |
  retainer
- |
  retaining
- |
  retainment
- |
  retake
- |
  retaken
- |
  retaliate
- |
  retaliation
- |
  retaliative
- |
  retaliator
- |
  retaliatory
- |
  retard
- |
  retardant
- |
  retardation
- |
  retarded
- |
  retarder
- |
  retaste
- |
  retaught
- |
  retch
- |
  reteach
- |
  retell
- |
  retelling
- |
  retention
- |
  retentive
- |
  retentively
- |
  retest
- |
  rethink
- |
  rethinking
- |
  rethought
- |
  reticence
- |
  reticent
- |
  reticently
- |
  reticulate
- |
  reticulated
- |
  reticulation
- |
  reticule
- |
  Reticulum
- |
  retie
- |
  retina
- |
  retinae
- |
  retinal
- |
  retinue
- |
  retire
- |
  retired
- |
  retiree
- |
  retirement
- |
  retiring
- |
  retiringness
- |
  retitle
- |
  retold
- |
  retook
- |
  retool
- |
  retort
- |
  retouch
- |
  retrace
- |
  retraceable
- |
  retract
- |
  retractable
- |
  retractible
- |
  retractile
- |
  retractility
- |
  retraction
- |
  retractive
- |
  retrain
- |
  retrainee
- |
  retraining
- |
  retranslate
- |
  retransmit
- |
  retread
- |
  retreat
- |
  retrench
- |
  retrenchment
- |
  retrial
- |
  retribution
- |
  retributive
- |
  retributory
- |
  retrievable
- |
  retrieval
- |
  retrieve
- |
  retriever
- |
  retro
- |
  retroaction
- |
  retroactive
- |
  retrocede
- |
  retrocession
- |
  retrod
- |
  retrodden
- |
  retrofire
- |
  retrofit
- |
  retrograde
- |
  retrogradely
- |
  retrogress
- |
  retronym
- |
  retrorocket
- |
  retrospect
- |
  retrousse
- |
  retrovirus
- |
  retry
- |
  retsina
- |
  retune
- |
  return
- |
  returnable
- |
  returnee
- |
  returner
- |
  returns
- |
  retype
- |
  Reuben
- |
  reunify
- |
  Reunion
- |
  reunion
- |
  reunite
- |
  reupholster
- |
  reusable
- |
  reuse
- |
  Reuther
- |
  revalidate
- |
  revalidation
- |
  revaluate
- |
  revaluation
- |
  revalue
- |
  revamp
- |
  revamped
- |
  revamping
- |
  revanche
- |
  revarnish
- |
  reveal
- |
  revealing
- |
  revealingly
- |
  reveille
- |
  revel
- |
  Revelation
- |
  revelation
- |
  Revelations
- |
  revelatory
- |
  reveler
- |
  reveller
- |
  revelry
- |
  revenant
- |
  revenge
- |
  revengeful
- |
  revenger
- |
  revenue
- |
  revenuer
- |
  reverb
- |
  reverberant
- |
  reverberate
- |
  reverberator
- |
  Revere
- |
  revere
- |
  revered
- |
  Reverence
- |
  reverence
- |
  Reverend
- |
  reverend
- |
  reverent
- |
  reverential
- |
  reverently
- |
  reverie
- |
  reverify
- |
  revers
- |
  reversal
- |
  reverse
- |
  reversely
- |
  reverser
- |
  reversible
- |
  reversibly
- |
  reversion
- |
  reversionary
- |
  revert
- |
  reverter
- |
  revertible
- |
  revery
- |
  revet
- |
  revetment
- |
  revetted
- |
  review
- |
  reviewer
- |
  revile
- |
  revilement
- |
  reviler
- |
  revisable
- |
  revisal
- |
  revise
- |
  reviser
- |
  revision
- |
  revisionism
- |
  revisionist
- |
  revisit
- |
  revisor
- |
  revisory
- |
  revitalise
- |
  revitalize
- |
  revivable
- |
  revival
- |
  revivalism
- |
  revivalist
- |
  revivalistic
- |
  revive
- |
  revived
- |
  reviver
- |
  revivify
- |
  revocable
- |
  revocation
- |
  revocatory
- |
  revokable
- |
  revoke
- |
  revoker
- |
  revolt
- |
  revolter
- |
  revolting
- |
  revoltingly
- |
  revolution
- |
  revolvable
- |
  revolve
- |
  revolver
- |
  revue
- |
  revulsion
- |
  revved
- |
  revving
- |
  rewaken
- |
  reward
- |
  rewarding
- |
  rewarm
- |
  rewash
- |
  reweave
- |
  rewed
- |
  reweigh
- |
  rewind
- |
  rewire
- |
  reword
- |
  rework
- |
  reworking
- |
  rewound
- |
  rewrap
- |
  rewrite
- |
  rewritten
- |
  rewrote
- |
  rewrought
- |
  Reykjavik
- |
  Reynold
- |
  Reynolds
- |
  rezone
- |
  Rhaetia
- |
  Rhaetian
- |
  rhapsodic
- |
  rhapsodical
- |
  rhapsodize
- |
  rhapsody
- |
  Rheims
- |
  Rhenish
- |
  rhenium
- |
  rheostat
- |
  rheostatic
- |
  rhesus
- |
  rhetoric
- |
  rhetorical
- |
  rhetorically
- |
  rhetorician
- |
  rheum
- |
  rheumatic
- |
  rheumatism
- |
  rheumatoid
- |
  rheumy
- |
  Rhine
- |
  Rhineland
- |
  Rhinelander
- |
  rhinestone
- |
  rhinestoned
- |
  rhinitis
- |
  rhino
- |
  rhinoceri
- |
  rhinoceros
- |
  rhizome
- |
  Rhoda
- |
  Rhodanus
- |
  Rhodes
- |
  Rhodesia
- |
  Rhodesian
- |
  rhodium
- |
  rhododendron
- |
  rhombi
- |
  rhomboid
- |
  rhomboidal
- |
  rhombus
- |
  Rhona
- |
  Rhone
- |
  rhubarb
- |
  rhyme
- |
  rhymer
- |
  rhymester
- |
  rhythm
- |
  rhythmic
- |
  rhythmical
- |
  rhythmically
- |
  rhythmless
- |
  ribald
- |
  ribaldry
- |
  riband
- |
  ribbed
- |
  ribber
- |
  ribbing
- |
  ribbon
- |
  ribbons
- |
  riboflavin
- |
  ribose
- |
  ribosomal
- |
  ribosome
- |
  Ricardo
- |
  ricer
- |
  Richard
- |
  Richardson
- |
  Richelieu
- |
  riches
- |
  richly
- |
  Richmond
- |
  richness
- |
  ricketiness
- |
  rickets
- |
  rickettsia
- |
  rickety
- |
  rickey
- |
  Rickover
- |
  rickrack
- |
  ricksha
- |
  rickshaw
- |
  ricochet
- |
  ricotta
- |
  ricrac
- |
  rictal
- |
  rictus
- |
  riddance
- |
  ridden
- |
  riddle
- |
  riddled
- |
  riddler
- |
  rider
- |
  riderless
- |
  ridership
- |
  ridge
- |
  ridgepole
- |
  ridgy
- |
  ridicule
- |
  ridiculous
- |
  ridiculously
- |
  riding
- |
  Riesling
- |
  rifely
- |
  rifeness
- |
  riffle
- |
  riffraff
- |
  rifle
- |
  rifleman
- |
  rifler
- |
  riflery
- |
  rifling
- |
  rifted
- |
  rifting
- |
  rigamarole
- |
  Rigel
- |
  rigger
- |
  rigging
- |
  Right
- |
  right
- |
  righteous
- |
  righteously
- |
  righter
- |
  rightful
- |
  rightfully
- |
  rightfulness
- |
  Rightism
- |
  rightism
- |
  rightist
- |
  rightly
- |
  rightmost
- |
  rightness
- |
  rights
- |
  rightsize
- |
  rightward
- |
  rigid
- |
  rigidity
- |
  rigidly
- |
  rigidness
- |
  rigmarole
- |
  rigor
- |
  rigorism
- |
  rigorist
- |
  rigorous
- |
  rigorously
- |
  rigorousness
- |
  rigors
- |
  rigour
- |
  Rilke
- |
  rille
- |
  rilled
- |
  Rimini
- |
  rimless
- |
  rimmed
- |
  ringer
- |
  ringgit
- |
  ringing
- |
  ringleader
- |
  ringlet
- |
  ringlike
- |
  ringmaster
- |
  ringside
- |
  ringworm
- |
  rinse
- |
  rinser
- |
  rioter
- |
  rioting
- |
  riotous
- |
  riotously
- |
  riotousness
- |
  riparian
- |
  ripcord
- |
  ripely
- |
  ripen
- |
  ripeness
- |
  ripoff
- |
  ripost
- |
  riposte
- |
  ripper
- |
  ripple
- |
  ripply
- |
  ripsaw
- |
  ripstop
- |
  riptide
- |
  risen
- |
  riser
- |
  risers
- |
  risibility
- |
  risible
- |
  risibly
- |
  rising
- |
  riskily
- |
  riskiness
- |
  risky
- |
  risotto
- |
  risque
- |
  ristra
- |
  ritard
- |
  ritual
- |
  ritualism
- |
  ritualist
- |
  ritualistic
- |
  ritualistize
- |
  ritualize
- |
  ritualized
- |
  ritually
- |
  rituals
- |
  ritzily
- |
  ritziness
- |
  ritzy
- |
  rival
- |
  rivalry
- |
  riven
- |
  river
- |
  Rivera
- |
  riverbank
- |
  riverbed
- |
  riverboat
- |
  riverfront
- |
  riverlike
- |
  Riverside
- |
  riverside
- |
  rivet
- |
  riveter
- |
  riveting
- |
  rivetingly
- |
  Riviera
- |
  rivulet
- |
  Riyadh
- |
  riyal
- |
  roach
- |
  roadbed
- |
  roadblock
- |
  roadhog
- |
  roadhouse
- |
  roadie
- |
  roadkill
- |
  roadrunner
- |
  roads
- |
  roadshow
- |
  roadside
- |
  roadstead
- |
  roadster
- |
  roadway
- |
  roadwork
- |
  roadworthy
- |
  roamer
- |
  Roanoke
- |
  roarer
- |
  roaring
- |
  roast
- |
  roaster
- |
  robber
- |
  robbery
- |
  Robbins
- |
  Robert
- |
  Roberta
- |
  Roberto
- |
  Robeson
- |
  Robespierre
- |
  Robin
- |
  robin
- |
  Robinson
- |
  robot
- |
  robotic
- |
  robotically
- |
  roboticist
- |
  robotics
- |
  robotize
- |
  robust
- |
  robustly
- |
  robustness
- |
  Robyn
- |
  rocaille
- |
  rocailles
- |
  Rochambeau
- |
  Rochelle
- |
  Rochester
- |
  rockabilly
- |
  rockbound
- |
  Rockefeller
- |
  rocker
- |
  rocket
- |
  rocketry
- |
  rockfall
- |
  rockfish
- |
  Rockford
- |
  Rockies
- |
  rockiness
- |
  Rockingham
- |
  rocklike
- |
  rocks
- |
  Rockville
- |
  Rockwell
- |
  Rocky
- |
  rocky
- |
  Rococo
- |
  rococo
- |
  rodent
- |
  rodeo
- |
  Roderick
- |
  Rodger
- |
  Rodgers
- |
  Rodin
- |
  Rodney
- |
  rodomontade
- |
  roebuck
- |
  Roentgen
- |
  roentgen
- |
  Roethke
- |
  Roger
- |
  roger
- |
  Rogers
- |
  Roget
- |
  rogue
- |
  roguery
- |
  roguish
- |
  roguishly
- |
  roguishness
- |
  roily
- |
  roister
- |
  roisterer
- |
  roisterous
- |
  Roland
- |
  Rolland
- |
  rollback
- |
  roller
- |
  Rollerblade
- |
  rollerskate
- |
  rollick
- |
  rollicking
- |
  Rollin
- |
  rolling
- |
  rollover
- |
  Rolvaag
- |
  Romagna
- |
  romaine
- |
  Roman
- |
  roman
- |
  Romance
- |
  romance
- |
  romancer
- |
  Romanesque
- |
  Romani
- |
  Romania
- |
  Romanian
- |
  Romanist
- |
  romanization
- |
  Romanize
- |
  romanize
- |
  Romano
- |
  Romanoff
- |
  Romanov
- |
  Romans
- |
  Romansch
- |
  Romansh
- |
  Romantic
- |
  romantic
- |
  romantically
- |
  Romanticism
- |
  romanticism
- |
  romanticist
- |
  romanticize
- |
  Romany
- |
  Romberg
- |
  Romblon
- |
  Romeo
- |
  Rommel
- |
  romper
- |
  rompers
- |
  Romulus
- |
  Ronal
- |
  Ronald
- |
  Ronda
- |
  ronde
- |
  rondeau
- |
  rondel
- |
  rondo
- |
  Ronnie
- |
  Ronny
- |
  Rontgen
- |
  roofed
- |
  roofer
- |
  roofie
- |
  roofing
- |
  roofless
- |
  rooftop
- |
  rooftree
- |
  rookery
- |
  rookie
- |
  roomer
- |
  roomette
- |
  roomful
- |
  roominess
- |
  roommate
- |
  rooms
- |
  roomy
- |
  Roosevelt
- |
  roost
- |
  rooster
- |
  rooted
- |
  rooter
- |
  rootless
- |
  rootlet
- |
  rootlike
- |
  roots
- |
  rootstock
- |
  ropes
- |
  Roquefort
- |
  rorqual
- |
  Rosalie
- |
  Rosalind
- |
  Rosalyn
- |
  Rosamond
- |
  Rosamund
- |
  Rosario
- |
  rosary
- |
  Roscoe
- |
  Roseanne
- |
  roseate
- |
  Roseau
- |
  rosebud
- |
  rosebush
- |
  Roselyn
- |
  Rosemarie
- |
  Rosemary
- |
  rosemary
- |
  Rosenberg
- |
  Rosetta
- |
  rosette
- |
  rosewater
- |
  rosewood
- |
  Rosicrucian
- |
  rosily
- |
  rosin
- |
  rosiness
- |
  rosiny
- |
  Rosita
- |
  Roslyn
- |
  Rossetti
- |
  Rossini
- |
  Rostand
- |
  roster
- |
  Rostock
- |
  Rostov
- |
  rostra
- |
  rostrate
- |
  rostrum
- |
  Roswell
- |
  rotary
- |
  rotatable
- |
  rotate
- |
  rotating
- |
  rotation
- |
  rotational
- |
  rotator
- |
  rotatory
- |
  rotgut
- |
  Rothko
- |
  Rothschild
- |
  rotisserie
- |
  rotogravure
- |
  rotor
- |
  rototill
- |
  rototiller
- |
  rotten
- |
  rottenness
- |
  rottenstone
- |
  Rotterdam
- |
  rottweiler
- |
  rotund
- |
  rotunda
- |
  rotundity
- |
  rotundly
- |
  rotundness
- |
  Rouault
- |
  rouble
- |
  Rouen
- |
  rouge
- |
  rough
- |
  roughage
- |
  roughen
- |
  rougher
- |
  roughhewn
- |
  roughhouse
- |
  roughly
- |
  roughneck
- |
  roughness
- |
  roughshod
- |
  roulade
- |
  roulette
- |
  Roumania
- |
  Roumanian
- |
  round
- |
  roundabout
- |
  rounded
- |
  roundel
- |
  roundelay
- |
  roundheel
- |
  roundhouse
- |
  roundish
- |
  roundly
- |
  roundness
- |
  rounds
- |
  roundtable
- |
  roundtrip
- |
  roundup
- |
  roundworm
- |
  rouse
- |
  rouser
- |
  rousing
- |
  Rousseau
- |
  roust
- |
  roustabout
- |
  route
- |
  routeman
- |
  router
- |
  routine
- |
  routinely
- |
  routinize
- |
  rover
- |
  roving
- |
  rowboat
- |
  rowdily
- |
  rowdiness
- |
  rowdy
- |
  rowdyish
- |
  rowdyism
- |
  rowel
- |
  Rowena
- |
  rower
- |
  rowing
- |
  Rowland
- |
  Roxanne
- |
  Royal
- |
  royal
- |
  royalist
- |
  royally
- |
  royalties
- |
  royalty
- |
  Royce
- |
  Ruanda
- |
  rubati
- |
  rubato
- |
  rubber
- |
  rubberiness
- |
  rubberize
- |
  rubberneck
- |
  rubbernecker
- |
  rubbery
- |
  rubbing
- |
  rubbish
- |
  rubbishy
- |
  rubble
- |
  rubbly
- |
  rubdown
- |
  rubel
- |
  rubella
- |
  Ruben
- |
  Rubenesque
- |
  Rubens
- |
  rubescent
- |
  Rubicon
- |
  rubicund
- |
  rubicundity
- |
  rubidium
- |
  rubiginous
- |
  Rubinstein
- |
  ruble
- |
  rubric
- |
  rubrical
- |
  rubricate
- |
  rubrication
- |
  rubricator
- |
  rucksack
- |
  ruckus
- |
  ruction
- |
  rudder
- |
  rudderless
- |
  ruddily
- |
  ruddiness
- |
  ruddy
- |
  rudely
- |
  rudeness
- |
  rudiment
- |
  rudimentary
- |
  rudiments
- |
  Rudolf
- |
  Rudolph
- |
  rueful
- |
  ruefully
- |
  ruefulness
- |
  rufescence
- |
  rufescent
- |
  ruffed
- |
  ruffian
- |
  ruffianly
- |
  ruffle
- |
  ruffled
- |
  ruffler
- |
  ruffly
- |
  rufiyaa
- |
  rufous
- |
  Rufus
- |
  Rugby
- |
  rugby
- |
  rugged
- |
  ruggedize
- |
  ruggedly
- |
  ruggedness
- |
  rugose
- |
  rugosity
- |
  ruinable
- |
  ruination
- |
  ruined
- |
  ruinous
- |
  ruinously
- |
  ruins
- |
  ruled
- |
  ruler
- |
  ruling
- |
  Rumania
- |
  Rumanian
- |
  rumba
- |
  rumble
- |
  rumbler
- |
  rumbling
- |
  rumblings
- |
  rumbly
- |
  rumbustious
- |
  rumen
- |
  rumina
- |
  ruminal
- |
  ruminant
- |
  ruminantly
- |
  ruminate
- |
  rumination
- |
  ruminative
- |
  ruminatively
- |
  ruminator
- |
  rummage
- |
  rummager
- |
  rummy
- |
  rumor
- |
  rumored
- |
  rumormonger
- |
  rumour
- |
  rumoured
- |
  rumple
- |
  rumpled
- |
  rumply
- |
  rumpus
- |
  rumrunner
- |
  runabout
- |
  runagate
- |
  runaround
- |
  runaway
- |
  rundown
- |
  runes
- |
  runic
- |
  runless
- |
  runlet
- |
  runnel
- |
  runner
- |
  running
- |
  runny
- |
  runoff
- |
  runtish
- |
  runty
- |
  runway
- |
  rupee
- |
  Rupert
- |
  rupiah
- |
  rupture
- |
  rural
- |
  ruralism
- |
  rurally
- |
  Rushdie
- |
  rushed
- |
  rusher
- |
  Rushmore
- |
  rushy
- |
  Ruskin
- |
  Ruskinian
- |
  Russel
- |
  Russell
- |
  russet
- |
  russety
- |
  Russia
- |
  Russian
- |
  Rustbelt
- |
  rustic
- |
  rustically
- |
  rusticate
- |
  rustication
- |
  rusticity
- |
  rustily
- |
  rustiness
- |
  rustle
- |
  rustler
- |
  rustling
- |
  rustproof
- |
  rusty
- |
  rutabaga
- |
  Rutgers
- |
  Ruthann
- |
  Ruthenia
- |
  Ruthenian
- |
  ruthenium
- |
  Rutherford
- |
  ruthless
- |
  ruthlessly
- |
  ruthlessness
- |
  rutting
- |
  rutty
- |
  Ruwenzori
- |
  Rwanda
- |
  Rwandan
- |
  Ryazan
- |
  Rybinsk
- |
  Ryukyu
- |
  Ryukyuan
- |
  Saarland
- |
  Sabah
- |
  Sabbath
- |
  sabbath
- |
  Sabbatical
- |
  sabbatical
- |
  saber
- |
  Sabin
- |
  Sabine
- |
  sable
- |
  sables
- |
  sabot
- |
  sabotage
- |
  saboteur
- |
  Sabra
- |
  sabra
- |
  sabre
- |
  Sacagawea
- |
  Sacajawea
- |
  saccharin
- |
  saccharine
- |
  Sacco
- |
  sacerdotal
- |
  sachem
- |
  sachet
- |
  Sachs
- |
  sackcloth
- |
  sacker
- |
  sackful
- |
  sacking
- |
  sacra
- |
  sacral
- |
  sacrality
- |
  Sacrament
- |
  sacrament
- |
  sacramental
- |
  Sacramento
- |
  sacraria
- |
  sacrarium
- |
  sacred
- |
  sacredly
- |
  sacredness
- |
  sacrifice
- |
  sacrificer
- |
  sacrificial
- |
  sacrilege
- |
  sacrilegious
- |
  sacrist
- |
  sacristan
- |
  sacristy
- |
  sacroiliac
- |
  sacrosanct
- |
  sacrosanctly
- |
  sacrum
- |
  Sadat
- |
  sadden
- |
  saddened
- |
  saddening
- |
  saddle
- |
  saddlebag
- |
  saddlebow
- |
  Sadducean
- |
  Sadducee
- |
  Sadie
- |
  sadiron
- |
  sadism
- |
  sadist
- |
  sadistic
- |
  sadistically
- |
  sadly
- |
  sadness
- |
  Safar
- |
  safari
- |
  safecracker
- |
  safecracking
- |
  safeguard
- |
  safekeeping
- |
  safelight
- |
  safely
- |
  safeness
- |
  safety
- |
  safflower
- |
  saffron
- |
  sagacious
- |
  sagaciously
- |
  sagacity
- |
  Sagamihara
- |
  sagamore
- |
  sagebrush
- |
  sagely
- |
  sageness
- |
  saggy
- |
  Saginaw
- |
  Sagitta
- |
  Sagittarian
- |
  Sagittarius
- |
  saguaro
- |
  Saguenay
- |
  Sahaptin
- |
  Sahara
- |
  Saharan
- |
  Saharian
- |
  Sahel
- |
  Sahelian
- |
  sahib
- |
  sahuaro
- |
  Saigon
- |
  sailboard
- |
  sailboarder
- |
  sailboarding
- |
  sailboat
- |
  sailcloth
- |
  sailfish
- |
  sailing
- |
  sailor
- |
  sailplane
- |
  saint
- |
  saintdom
- |
  sainted
- |
  sainthood
- |
  saintlike
- |
  saintliness
- |
  saintly
- |
  Saipan
- |
  Saipanese
- |
  saith
- |
  Sakai
- |
  Sakhalin
- |
  Sakharov
- |
  salaam
- |
  salability
- |
  salable
- |
  salacious
- |
  salaciously
- |
  salacity
- |
  salad
- |
  Saladin
- |
  Salamanca
- |
  salamander
- |
  salami
- |
  Salamis
- |
  salaried
- |
  salary
- |
  Salazar
- |
  saleable
- |
  Salem
- |
  Salerno
- |
  sales
- |
  salesclerk
- |
  salesgirl
- |
  saleslady
- |
  salesman
- |
  salesmanship
- |
  salespeople
- |
  salesperson
- |
  saleswoman
- |
  Salford
- |
  salience
- |
  saliency
- |
  salient
- |
  saliently
- |
  Salinas
- |
  saline
- |
  Salinger
- |
  salinity
- |
  salinization
- |
  salinize
- |
  Salisbury
- |
  Salish
- |
  Salishan
- |
  saliva
- |
  salivary
- |
  salivate
- |
  salivation
- |
  Sallie
- |
  sallow
- |
  sallowish
- |
  sallowly
- |
  sallowness
- |
  Sallust
- |
  Sally
- |
  sally
- |
  salmagundi
- |
  salmon
- |
  salmonella
- |
  salmonellae
- |
  Salome
- |
  Salon
- |
  salon
- |
  Salonika
- |
  saloon
- |
  Salop
- |
  salsa
- |
  saltation
- |
  saltatory
- |
  saltcellar
- |
  salted
- |
  Saltillo
- |
  saltily
- |
  saltine
- |
  saltiness
- |
  saltpeter
- |
  saltpetre
- |
  salts
- |
  saltshaker
- |
  saltwater
- |
  salty
- |
  salubrious
- |
  salubriously
- |
  salubrity
- |
  salutarily
- |
  salutariness
- |
  salutary
- |
  salutation
- |
  salutational
- |
  salutatorian
- |
  salutatory
- |
  salute
- |
  Salvador
- |
  Salvadoran
- |
  Salvadorean
- |
  Salvadorian
- |
  salvage
- |
  salvageable
- |
  salvager
- |
  salvation
- |
  salvational
- |
  Salvatore
- |
  salve
- |
  salver
- |
  salvia
- |
  salvo
- |
  Salween
- |
  Salzburg
- |
  Samantha
- |
  Samar
- |
  Samara
- |
  Samaria
- |
  Samarinda
- |
  Samaritan
- |
  samaritan
- |
  samarium
- |
  Samarkand
- |
  Samarqand
- |
  samba
- |
  sameness
- |
  Samian
- |
  samizdat
- |
  Sammie
- |
  Sammy
- |
  Samnite
- |
  Samnium
- |
  Samoa
- |
  Samoan
- |
  Samos
- |
  Samoset
- |
  samovar
- |
  Samoyed
- |
  sampan
- |
  sample
- |
  sampler
- |
  sampling
- |
  samsara
- |
  samsaric
- |
  Samson
- |
  Samsun
- |
  Samuel
- |
  samurai
- |
  Sanaa
- |
  sanative
- |
  sanatoria
- |
  sanatorium
- |
  Sanchung
- |
  sancta
- |
  sanctifier
- |
  sanctify
- |
  sanctimony
- |
  sanction
- |
  sanctionable
- |
  sanctions
- |
  sanctity
- |
  sanctuary
- |
  sanctum
- |
  sandal
- |
  sandaled
- |
  sandalwood
- |
  sandbag
- |
  sandbank
- |
  sandbar
- |
  sandblast
- |
  sandblaster
- |
  sandbox
- |
  Sandburg
- |
  sandcastle
- |
  sander
- |
  sandhog
- |
  sandiness
- |
  sandlot
- |
  sandlotter
- |
  sandman
- |
  sandpaper
- |
  sandpiper
- |
  Sandra
- |
  sandstone
- |
  sandstorm
- |
  Sandwich
- |
  sandwich
- |
  Sandy
- |
  sandy
- |
  sanely
- |
  saneness
- |
  Sanford
- |
  Sanforized
- |
  Sanger
- |
  sangfroid
- |
  sangria
- |
  sanguinarily
- |
  sanguinary
- |
  sanguine
- |
  sanguinely
- |
  sanguineness
- |
  sanguineous
- |
  sanguinity
- |
  sanitaria
- |
  sanitarian
- |
  sanitarily
- |
  sanitarium
- |
  sanitary
- |
  sanitation
- |
  sanitize
- |
  sanity
- |
  Sanscrit
- |
  sansei
- |
  Sanskrit
- |
  Sanskritist
- |
  Santa
- |
  Santayana
- |
  Santee
- |
  Santeria
- |
  Santiago
- |
  Saone
- |
  Saphar
- |
  sapid
- |
  sapidity
- |
  sapience
- |
  sapient
- |
  sapiently
- |
  sapless
- |
  sapling
- |
  sapodilla
- |
  saponaceous
- |
  saponifiable
- |
  saponified
- |
  saponify
- |
  sapper
- |
  Sapphic
- |
  sapphic
- |
  sapphics
- |
  sapphire
- |
  sapphism
- |
  Sappho
- |
  sappiness
- |
  Sapporo
- |
  sappy
- |
  saprophyte
- |
  saprophytic
- |
  sapsucker
- |
  sapwood
- |
  Saracen
- |
  Saragossa
- |
  Sarah
- |
  Sarajevo
- |
  Saralee
- |
  saran
- |
  sarape
- |
  Sarasota
- |
  Saratoga
- |
  Saratov
- |
  Sarawak
- |
  sarcasm
- |
  sarcastic
- |
  sarcoid
- |
  sarcoma
- |
  sarcomata
- |
  sarcophagi
- |
  sarcophagus
- |
  sardine
- |
  Sardinia
- |
  Sardinian
- |
  Sardis
- |
  sardonic
- |
  sardonically
- |
  sardonicism
- |
  saree
- |
  sargasso
- |
  sarge
- |
  Sargent
- |
  Sargon
- |
  Sarmatia
- |
  Sarmatian
- |
  sarong
- |
  Saroyan
- |
  sarsaparilla
- |
  sartorial
- |
  sartorially
- |
  Sartre
- |
  sashay
- |
  Saskatchewan
- |
  Saskatoon
- |
  Sasquatch
- |
  sassafras
- |
  sassily
- |
  sassiness
- |
  sassy
- |
  Satan
- |
  satang
- |
  satanic
- |
  satanical
- |
  satanically
- |
  Satanism
- |
  satanism
- |
  Satanist
- |
  satanist
- |
  satanistic
- |
  satchel
- |
  sateen
- |
  sateless
- |
  satellite
- |
  satiable
- |
  satiate
- |
  satiation
- |
  satiety
- |
  satin
- |
  satinwood
- |
  satiny
- |
  satire
- |
  satiric
- |
  satirical
- |
  satirically
- |
  satirist
- |
  satirization
- |
  satirize
- |
  satisfaction
- |
  satisfactory
- |
  satisfied
- |
  satisfy
- |
  satisfying
- |
  satisfyingly
- |
  satori
- |
  satrap
- |
  saturable
- |
  saturate
- |
  saturated
- |
  saturates
- |
  saturation
- |
  Saturday
- |
  Saturn
- |
  Saturnalia
- |
  saturnalia
- |
  saturnalian
- |
  saturnine
- |
  saturninely
- |
  satyagraha
- |
  Satyr
- |
  satyr
- |
  satyriasis
- |
  satyric
- |
  sauce
- |
  saucepan
- |
  saucer
- |
  saucily
- |
  sauciness
- |
  saucy
- |
  saudade
- |
  Saudi
- |
  sauerbraten
- |
  sauerkraut
- |
  sauna
- |
  Saundra
- |
  saunter
- |
  saunterer
- |
  saurian
- |
  sauropod
- |
  sausage
- |
  Saussure
- |
  saute
- |
  sauterne
- |
  Sauternes
- |
  sauternes
- |
  savable
- |
  savage
- |
  savagely
- |
  savageness
- |
  savagery
- |
  Savaii
- |
  savanna
- |
  Savannah
- |
  savannah
- |
  savant
- |
  saveable
- |
  saver
- |
  saving
- |
  savings
- |
  Savior
- |
  savior
- |
  saviour
- |
  Savonarola
- |
  savor
- |
  savorer
- |
  savorily
- |
  savoriness
- |
  savorless
- |
  savory
- |
  savour
- |
  savoury
- |
  Savoy
- |
  Savoyard
- |
  savvy
- |
  sawbuck
- |
  sawdust
- |
  sawer
- |
  sawfish
- |
  sawfly
- |
  sawhorse
- |
  sawmill
- |
  sawyer
- |
  saxifrage
- |
  Saxon
- |
  Saxony
- |
  saxophone
- |
  saxophonist
- |
  sayer
- |
  Sayers
- |
  saying
- |
  sayonara
- |
  scabbard
- |
  scabbed
- |
  scabbiness
- |
  scabby
- |
  scabies
- |
  scabietic
- |
  scablands
- |
  scablike
- |
  scabrous
- |
  scabrously
- |
  scabrousness
- |
  scads
- |
  scaffold
- |
  scaffolding
- |
  scalable
- |
  scalar
- |
  scalawag
- |
  scald
- |
  scalding
- |
  Scaldis
- |
  scale
- |
  scaled
- |
  scaleless
- |
  scalene
- |
  scalepan
- |
  scales
- |
  Scalia
- |
  scaliness
- |
  scallion
- |
  scallop
- |
  scalloped
- |
  scalloper
- |
  scalloping
- |
  scallywag
- |
  scalp
- |
  scalpel
- |
  scalper
- |
  scaly
- |
  scamp
- |
  scamper
- |
  scamperer
- |
  scampi
- |
  scandal
- |
  scandalize
- |
  scandalizer
- |
  scandalous
- |
  scandalously
- |
  scandent
- |
  Scandinavia
- |
  Scandinavian
- |
  scandium
- |
  scannable
- |
  scanner
- |
  scanning
- |
  scansion
- |
  scant
- |
  scantily
- |
  scantiness
- |
  scantling
- |
  scantly
- |
  scantness
- |
  scanty
- |
  scapegoat
- |
  scapegoater
- |
  scapegoating
- |
  scapegoatism
- |
  scapegrace
- |
  scapula
- |
  scapulae
- |
  scapular
- |
  scarab
- |
  scaramouch
- |
  Scarborough
- |
  scarce
- |
  scarcely
- |
  scarceness
- |
  scarcity
- |
  scare
- |
  scarecrow
- |
  scared
- |
  scarf
- |
  scarify
- |
  scarifying
- |
  scarily
- |
  scariness
- |
  scarlatina
- |
  Scarlatti
- |
  scarlet
- |
  scarp
- |
  scarves
- |
  scary
- |
  scathe
- |
  scathing
- |
  scathingly
- |
  scatologic
- |
  scatological
- |
  scatology
- |
  scatter
- |
  scatterbrain
- |
  scattered
- |
  scatterer
- |
  scattering
- |
  scattershot
- |
  scavenge
- |
  scavenger
- |
  scenario
- |
  scenarist
- |
  scene
- |
  scenery
- |
  scenic
- |
  scenically
- |
  scenographer
- |
  scenography
- |
  scent
- |
  scented
- |
  scentless
- |
  scepter
- |
  sceptered
- |
  sceptic
- |
  sceptical
- |
  sceptically
- |
  scepticism
- |
  sceptre
- |
  Scheat
- |
  Schedar
- |
  schedule
- |
  scheduler
- |
  Scheherazade
- |
  Schelde
- |
  Scheldt
- |
  Schelling
- |
  schema
- |
  schemata
- |
  schematic
- |
  schematize
- |
  scheme
- |
  schemer
- |
  scheming
- |
  Schenectady
- |
  scherzi
- |
  scherzo
- |
  Schiller
- |
  schilling
- |
  schism
- |
  schismatic
- |
  schist
- |
  schistose
- |
  schizo
- |
  schizoid
- |
  schlemiel
- |
  schlep
- |
  schlepp
- |
  schlepper
- |
  Schleswig
- |
  Schliemann
- |
  schlock
- |
  schlocky
- |
  schmaltz
- |
  schmaltzy
- |
  schmalz
- |
  schmear
- |
  schmeer
- |
  Schmidt
- |
  schmo
- |
  schmoe
- |
  schmooze
- |
  schmuck
- |
  schnapps
- |
  schnaps
- |
  schnauzer
- |
  schnitzel
- |
  schnook
- |
  schnorrer
- |
  schnoz
- |
  schnozzle
- |
  scholar
- |
  scholarly
- |
  scholarship
- |
  scholastic
- |
  Schonberg
- |
  school
- |
  schoolbook
- |
  schoolboy
- |
  schoolchild
- |
  schooled
- |
  schoolfellow
- |
  schoolgirl
- |
  schoolhouse
- |
  schooling
- |
  schoolmarm
- |
  schoolmaster
- |
  schoolmate
- |
  schoolroom
- |
  schoolwork
- |
  schoolyard
- |
  schooner
- |
  Schopenhauer
- |
  schrod
- |
  Schrodinger
- |
  Schubert
- |
  Schulz
- |
  Schumann
- |
  schuss
- |
  schussboomer
- |
  schwa
- |
  Schweitzer
- |
  sciatic
- |
  sciatica
- |
  sciatically
- |
  science
- |
  scientific
- |
  scientist
- |
  scilicet
- |
  Scilly
- |
  scimitar
- |
  scintilla
- |
  scintillant
- |
  scintillate
- |
  sciolism
- |
  sciolist
- |
  sciolistic
- |
  scion
- |
  Scipio
- |
  scirocco
- |
  scission
- |
  scissor
- |
  scissors
- |
  sclera
- |
  scleral
- |
  scleroses
- |
  sclerosis
- |
  sclerotic
- |
  scoff
- |
  scoffer
- |
  scofflaw
- |
  scold
- |
  scolder
- |
  scolding
- |
  scoliosis
- |
  scoliotic
- |
  sconce
- |
  scone
- |
  scoop
- |
  scooper
- |
  scoot
- |
  scooter
- |
  scope
- |
  Scopes
- |
  scorbutic
- |
  scorbutical
- |
  scorch
- |
  scorched
- |
  scorcher
- |
  scorching
- |
  score
- |
  scoreboard
- |
  scorecard
- |
  scorekeeper
- |
  scoreless
- |
  scorer
- |
  scores
- |
  scoria
- |
  scoriaceous
- |
  scoriae
- |
  scorn
- |
  scorner
- |
  scornful
- |
  scornfully
- |
  scornfulness
- |
  Scorpio
- |
  scorpion
- |
  Scorpius
- |
  Scotch
- |
  scotch
- |
  Scotchman
- |
  Scotchwoman
- |
  Scotia
- |
  Scotland
- |
  scotopic
- |
  Scots
- |
  Scotsman
- |
  Scotswoman
- |
  Scott
- |
  Scottie
- |
  Scottish
- |
  Scottsdale
- |
  Scotty
- |
  scoundrel
- |
  scoundrelly
- |
  scour
- |
  scourer
- |
  scourge
- |
  scourger
- |
  scours
- |
  Scout
- |
  scout
- |
  scouting
- |
  scoutmaster
- |
  scowl
- |
  scowler
- |
  scowlingly
- |
  Scrabble
- |
  scrabble
- |
  scrabbler
- |
  scragginess
- |
  scraggly
- |
  scraggy
- |
  scram
- |
  scramble
- |
  scrambled
- |
  scrambler
- |
  Scranton
- |
  scrap
- |
  scrapbook
- |
  scrape
- |
  scraper
- |
  scrapheap
- |
  scraping
- |
  scrapper
- |
  scrappily
- |
  scrappiness
- |
  scrappy
- |
  scraps
- |
  scrapyard
- |
  scratch
- |
  scratcher
- |
  scratchily
- |
  scratchiness
- |
  scratchy
- |
  scrawl
- |
  scrawly
- |
  scrawniness
- |
  scrawny
- |
  scream
- |
  screamer
- |
  screaming
- |
  scree
- |
  screech
- |
  screechy
- |
  screed
- |
  screen
- |
  screener
- |
  screening
- |
  screenplay
- |
  screenwriter
- |
  screw
- |
  screwball
- |
  screwdriver
- |
  screwiness
- |
  screwworm
- |
  screwy
- |
  scribal
- |
  scribble
- |
  scribbler
- |
  scribbles
- |
  Scribe
- |
  scribe
- |
  scriber
- |
  scrim
- |
  scrimmage
- |
  scrimmager
- |
  scrimp
- |
  scrimper
- |
  scrimshander
- |
  scrimshaw
- |
  scrip
- |
  script
- |
  scripted
- |
  scriptoria
- |
  scriptorium
- |
  Scriptural
- |
  scriptural
- |
  scripturally
- |
  Scripture
- |
  scripture
- |
  Scriptures
- |
  scriptwriter
- |
  scrivener
- |
  scrod
- |
  scrofula
- |
  scrofulous
- |
  scroll
- |
  Scrooge
- |
  scrooge
- |
  scrota
- |
  scrotal
- |
  scrotum
- |
  scrounge
- |
  scrounger
- |
  scrounginess
- |
  scroungy
- |
  scrub
- |
  scrubber
- |
  scrubby
- |
  scrubwoman
- |
  scruff
- |
  scruffily
- |
  scruffiness
- |
  scruffy
- |
  scrum
- |
  scrumptious
- |
  scrunch
- |
  scrunchie
- |
  scrunchy
- |
  scruple
- |
  scruples
- |
  scrupulosity
- |
  scrupulous
- |
  scrupulously
- |
  scrutinise
- |
  scrutinize
- |
  scrutinizer
- |
  scrutiny
- |
  scuba
- |
  scuff
- |
  scuffle
- |
  scuffler
- |
  scull
- |
  sculler
- |
  scullery
- |
  scullion
- |
  sculls
- |
  sculpt
- |
  Sculptor
- |
  sculptor
- |
  sculptress
- |
  sculptural
- |
  sculpture
- |
  sculptured
- |
  scumbag
- |
  scumble
- |
  scummy
- |
  scupper
- |
  scuppers
- |
  scurf
- |
  scurfiness
- |
  scurfy
- |
  scurrility
- |
  scurrilous
- |
  scurrilously
- |
  scurry
- |
  scurvily
- |
  scurviness
- |
  scurvy
- |
  scutage
- |
  scutcheon
- |
  scuttle
- |
  scuttlebutt
- |
  Scutum
- |
  scuzzy
- |
  Scylla
- |
  scythe
- |
  Scythia
- |
  Scythian
- |
  seabed
- |
  seabird
- |
  seaboard
- |
  seaborgium
- |
  seacoast
- |
  seafarer
- |
  seafaring
- |
  seafood
- |
  seagoing
- |
  seagull
- |
  seahorse
- |
  sealable
- |
  sealane
- |
  sealant
- |
  sealed
- |
  sealer
- |
  sealskin
- |
  Seaman
- |
  seaman
- |
  seamanship
- |
  seaminess
- |
  seamless
- |
  seamlessly
- |
  seamount
- |
  seamstress
- |
  seamy
- |
  seance
- |
  seaplane
- |
  seaport
- |
  seaquake
- |
  search
- |
  searcher
- |
  searching
- |
  searchingly
- |
  searchlight
- |
  searing
- |
  seascape
- |
  seashell
- |
  seashore
- |
  seasick
- |
  seasickness
- |
  seaside
- |
  season
- |
  seasonable
- |
  seasonably
- |
  seasonal
- |
  seasonally
- |
  seasoned
- |
  seasoner
- |
  seasoning
- |
  seatbelt
- |
  seating
- |
  Seattle
- |
  seawall
- |
  seaward
- |
  seawards
- |
  seawater
- |
  seaway
- |
  seaweed
- |
  seaworthy
- |
  sebaceous
- |
  Sebastian
- |
  seborrhea
- |
  seborrheic
- |
  seborrhoea
- |
  secant
- |
  secco
- |
  secede
- |
  Secession
- |
  secession
- |
  secessional
- |
  secessionism
- |
  secessionist
- |
  seclude
- |
  secluded
- |
  seclusion
- |
  seclusive
- |
  second
- |
  secondarily
- |
  secondary
- |
  seconder
- |
  secondhand
- |
  secondly
- |
  seconds
- |
  secrecy
- |
  secret
- |
  secretarial
- |
  secretariat
- |
  secretary
- |
  secrete
- |
  secretion
- |
  secretionary
- |
  secretive
- |
  secretively
- |
  secretly
- |
  secretor
- |
  secretory
- |
  sectarian
- |
  sectarianism
- |
  sectarianize
- |
  sectary
- |
  section
- |
  sectional
- |
  sectionalism
- |
  sectionalist
- |
  sectionally
- |
  sector
- |
  sectoral
- |
  sectorial
- |
  secular
- |
  secularism
- |
  secularist
- |
  secularistic
- |
  secularity
- |
  secularize
- |
  secularizer
- |
  secularly
- |
  secure
- |
  securely
- |
  securement
- |
  securities
- |
  security
- |
  sedan
- |
  sedate
- |
  sedated
- |
  sedately
- |
  sedateness
- |
  sedation
- |
  sedative
- |
  sedentarily
- |
  sedentary
- |
  Seder
- |
  sedge
- |
  sedgy
- |
  sediment
- |
  sedimentary
- |
  sedimented
- |
  sedition
- |
  seditionist
- |
  seditious
- |
  seditiously
- |
  seduce
- |
  seducer
- |
  seducible
- |
  seduction
- |
  seductive
- |
  seductively
- |
  seductress
- |
  sedulity
- |
  sedulous
- |
  sedulously
- |
  sedulousness
- |
  sedum
- |
  seedbed
- |
  seedcase
- |
  seeder
- |
  seedily
- |
  seediness
- |
  seedless
- |
  seedlessness
- |
  seedling
- |
  seedpod
- |
  seedtime
- |
  seedy
- |
  seeing
- |
  seeker
- |
  seeming
- |
  seemingly
- |
  seemliness
- |
  seemly
- |
  seepage
- |
  seeress
- |
  seersucker
- |
  seesaw
- |
  seethe
- |
  seething
- |
  segment
- |
  segmental
- |
  segmentalize
- |
  segmentally
- |
  segmentation
- |
  segmented
- |
  Segovia
- |
  segregable
- |
  segregate
- |
  segregated
- |
  segregation
- |
  segregative
- |
  segregator
- |
  segue
- |
  seicento
- |
  seigneur
- |
  seigneurial
- |
  seignior
- |
  seigniorial
- |
  seignorial
- |
  Seine
- |
  seine
- |
  seiner
- |
  seismic
- |
  seismical
- |
  seismically
- |
  seismicity
- |
  seismogram
- |
  seismograph
- |
  seismography
- |
  seismologic
- |
  seismologist
- |
  seismology
- |
  seismometer
- |
  seitan
- |
  seizable
- |
  seize
- |
  seizer
- |
  seizure
- |
  seldom
- |
  seldomness
- |
  select
- |
  selectee
- |
  selection
- |
  selective
- |
  selectively
- |
  selectivity
- |
  selectman
- |
  selectness
- |
  selector
- |
  selectwoman
- |
  selenite
- |
  selenium
- |
  selenography
- |
  Seleucia
- |
  Seleucid
- |
  Seleucus
- |
  selfish
- |
  selfishly
- |
  selfishness
- |
  selfless
- |
  selflessly
- |
  selflessness
- |
  selfsame
- |
  Seljuk
- |
  Selkirk
- |
  seller
- |
  selloff
- |
  sellout
- |
  Selma
- |
  seltzer
- |
  selvage
- |
  selvaged
- |
  selvedge
- |
  selves
- |
  semantic
- |
  semantical
- |
  semantically
- |
  semantician
- |
  semanticist
- |
  semantics
- |
  semaphore
- |
  Semarang
- |
  semasiology
- |
  semblable
- |
  semblance
- |
  semen
- |
  semester
- |
  semiannual
- |
  semiannually
- |
  semiarid
- |
  semicircle
- |
  semicircular
- |
  semicolon
- |
  semidarkness
- |
  semidivine
- |
  semifinal
- |
  semifinalist
- |
  semiformal
- |
  semigloss
- |
  semiliquid
- |
  semiliterate
- |
  semilunar
- |
  semimonthly
- |
  seminal
- |
  seminally
- |
  seminar
- |
  seminarian
- |
  seminarist
- |
  seminary
- |
  Seminole
- |
  semiofficial
- |
  semiological
- |
  semiologist
- |
  semiology
- |
  semiotic
- |
  semiotically
- |
  semiotician
- |
  semioticism
- |
  semiotics
- |
  semiprecious
- |
  semiprivate
- |
  semipro
- |
  semiretired
- |
  semiskilled
- |
  semisoft
- |
  semisolid
- |
  semisweet
- |
  Semite
- |
  Semitic
- |
  Semitism
- |
  semitone
- |
  semitonic
- |
  semitrailer
- |
  semitropical
- |
  semivowel
- |
  semiweekly
- |
  semiyearly
- |
  semolina
- |
  sempiternal
- |
  sempiternity
- |
  sempstress
- |
  Semtex
- |
  Senate
- |
  senate
- |
  Senator
- |
  senator
- |
  senatorial
- |
  Sendai
- |
  sender
- |
  sendoff
- |
  Seneca
- |
  Senegal
- |
  Senegalese
- |
  senescence
- |
  senescent
- |
  senile
- |
  senilely
- |
  senility
- |
  Senior
- |
  senior
- |
  seniority
- |
  seniti
- |
  senna
- |
  Sennacherib
- |
  senor
- |
  senora
- |
  senores
- |
  senorita
- |
  sensate
- |
  sensation
- |
  sensational
- |
  sense
- |
  senseless
- |
  senselessly
- |
  senses
- |
  sensibility
- |
  sensible
- |
  sensibleness
- |
  sensibly
- |
  sensitive
- |
  sensitively
- |
  sensitivity
- |
  sensitize
- |
  sensor
- |
  sensoria
- |
  sensorium
- |
  sensory
- |
  sensual
- |
  sensualism
- |
  sensualist
- |
  sensuality
- |
  sensualize
- |
  sensually
- |
  sensualness
- |
  sensuosity
- |
  sensuous
- |
  sensuously
- |
  sensuousness
- |
  sente
- |
  sentence
- |
  sentential
- |
  sententially
- |
  sententious
- |
  sentience
- |
  sentiency
- |
  sentient
- |
  sentiently
- |
  sentiment
- |
  sentimental
- |
  sentimo
- |
  sentinel
- |
  sentry
- |
  Seoul
- |
  sepal
- |
  sepaled
- |
  sepalous
- |
  separability
- |
  separable
- |
  separably
- |
  separate
- |
  separated
- |
  separately
- |
  separateness
- |
  separates
- |
  separation
- |
  separatism
- |
  separatist
- |
  separative
- |
  separator
- |
  Sephardi
- |
  Sephardic
- |
  sepia
- |
  seppuku
- |
  sepses
- |
  sepsis
- |
  septa
- |
  September
- |
  septennial
- |
  septennially
- |
  septet
- |
  septette
- |
  septic
- |
  septically
- |
  septicemia
- |
  septicemic
- |
  septicity
- |
  septillion
- |
  septillionth
- |
  Septuagint
- |
  septum
- |
  septuplet
- |
  sepulcher
- |
  sepulchral
- |
  sepulchrally
- |
  sepulchre
- |
  sepulture
- |
  sequacious
- |
  sequaciously
- |
  sequacity
- |
  sequel
- |
  sequela
- |
  sequelae
- |
  sequence
- |
  sequencing
- |
  sequent
- |
  sequential
- |
  sequentially
- |
  sequently
- |
  sequester
- |
  sequestrable
- |
  sequestrate
- |
  sequestrated
- |
  sequestrator
- |
  sequin
- |
  sequined
- |
  sequinned
- |
  sequoia
- |
  Sequoya
- |
  Sequoyah
- |
  Seraglio
- |
  seraglio
- |
  serape
- |
  seraph
- |
  seraphic
- |
  seraphical
- |
  seraphically
- |
  seraphim
- |
  Serbia
- |
  Serbian
- |
  serenade
- |
  serenader
- |
  serendipity
- |
  Serene
- |
  serene
- |
  serenely
- |
  sereneness
- |
  Serengeti
- |
  serenity
- |
  serfage
- |
  serfdom
- |
  serge
- |
  Sergeant
- |
  sergeant
- |
  serial
- |
  serialism
- |
  serialist
- |
  seriality
- |
  serialize
- |
  serially
- |
  serials
- |
  seriatim
- |
  sericultural
- |
  sericulture
- |
  series
- |
  serif
- |
  seriffed
- |
  serigraph
- |
  serigrapher
- |
  serigraphy
- |
  seriocomic
- |
  serious
- |
  seriously
- |
  seriousness
- |
  sermon
- |
  sermonize
- |
  sermonizer
- |
  serologic
- |
  serological
- |
  serologist
- |
  serology
- |
  seronegative
- |
  seropositive
- |
  serotonin
- |
  serous
- |
  Serpens
- |
  serpent
- |
  serpentine
- |
  Serra
- |
  serrate
- |
  serrated
- |
  serration
- |
  serried
- |
  serum
- |
  servant
- |
  serve
- |
  server
- |
  service
- |
  serviceable
- |
  serviceably
- |
  serviceman
- |
  servicewoman
- |
  servile
- |
  servilely
- |
  servileness
- |
  servility
- |
  serving
- |
  servitor
- |
  servitude
- |
  servo
- |
  servomotor
- |
  sesame
- |
  sessile
- |
  session
- |
  sestet
- |
  sestina
- |
  setaceous
- |
  setaceously
- |
  setback
- |
  Seton
- |
  setscrew
- |
  settee
- |
  setter
- |
  setting
- |
  settle
- |
  settled
- |
  settlement
- |
  settler
- |
  settlor
- |
  setup
- |
  setups
- |
  Seurat
- |
  Seuss
- |
  Sevastopol
- |
  seven
- |
  seventeen
- |
  seventeenth
- |
  seventh
- |
  seventieth
- |
  seventy
- |
  sever
- |
  several
- |
  severally
- |
  severalty
- |
  severance
- |
  severe
- |
  severely
- |
  severeness
- |
  severity
- |
  Severn
- |
  Severus
- |
  Seville
- |
  Sevillian
- |
  sewage
- |
  Seward
- |
  sewer
- |
  sewerage
- |
  sewing
- |
  sexagenarian
- |
  sexagesimal
- |
  sexed
- |
  sexily
- |
  sexiness
- |
  sexism
- |
  sexist
- |
  sexless
- |
  sexlessly
- |
  sexlessness
- |
  sexological
- |
  sexologist
- |
  sexology
- |
  sexpot
- |
  Sextans
- |
  sextant
- |
  sextet
- |
  sextette
- |
  sextillion
- |
  sextillionth
- |
  Sexton
- |
  sexton
- |
  sextuple
- |
  sextuplet
- |
  sextuply
- |
  sexual
- |
  sexuality
- |
  sexually
- |
  Seychelles
- |
  Seymour
- |
  Sezession
- |
  sforzandi
- |
  sforzando
- |
  sforzati
- |
  sforzato
- |
  sgraffiti
- |
  sgraffito
- |
  Shaaban
- |
  Shabbat
- |
  shabbily
- |
  shabbiness
- |
  shabby
- |
  shack
- |
  shackle
- |
  shackles
- |
  shade
- |
  shaded
- |
  shades
- |
  shadily
- |
  shadiness
- |
  shading
- |
  shadow
- |
  shadowbox
- |
  shadowboxing
- |
  shadower
- |
  shadowiness
- |
  shadowy
- |
  shady
- |
  shaft
- |
  shagginess
- |
  shaggy
- |
  shaikh
- |
  shakable
- |
  shake
- |
  shakedown
- |
  shaken
- |
  shakeout
- |
  Shaker
- |
  shaker
- |
  Shakerism
- |
  Shakespeare
- |
  shakeup
- |
  shakily
- |
  shakiness
- |
  shako
- |
  shaky
- |
  shale
- |
  shaley
- |
  shall
- |
  shallop
- |
  shallot
- |
  shallow
- |
  shallowly
- |
  shallowness
- |
  shallows
- |
  shalom
- |
  shalt
- |
  shaman
- |
  shamanic
- |
  shamanism
- |
  shamanist
- |
  shamanistic
- |
  shamanize
- |
  shamble
- |
  shambles
- |
  shambling
- |
  shame
- |
  shamefaced
- |
  shamefacedly
- |
  shameful
- |
  shamefully
- |
  shamefulness
- |
  shameless
- |
  shamelessly
- |
  shammer
- |
  shammy
- |
  shampoo
- |
  shampooer
- |
  shamrock
- |
  Shandong
- |
  Shane
- |
  Shanghai
- |
  shanghai
- |
  shank
- |
  Shankar
- |
  Shannon
- |
  Shantung
- |
  shantung
- |
  shanty
- |
  shape
- |
  shaped
- |
  shapeless
- |
  shapelessly
- |
  shapeliness
- |
  shapely
- |
  shaper
- |
  shard
- |
  share
- |
  sharecrop
- |
  sharecropper
- |
  shareholder
- |
  shareholding
- |
  sharer
- |
  shareware
- |
  Shari
- |
  shark
- |
  sharkskin
- |
  Sharlene
- |
  Sharon
- |
  sharp
- |
  sharpen
- |
  sharpener
- |
  sharper
- |
  sharpie
- |
  sharply
- |
  sharpness
- |
  sharpshooter
- |
  sharpy
- |
  Sharron
- |
  Shasta
- |
  shatter
- |
  shattered
- |
  shattering
- |
  shatterproof
- |
  shave
- |
  shaven
- |
  shaver
- |
  shaves
- |
  Shavian
- |
  shaving
- |
  shavings
- |
  shawl
- |
  Shawn
- |
  Shawnee
- |
  Shawwal
- |
  shaykh
- |
  Shays
- |
  sheaf
- |
  shear
- |
  shearer
- |
  shearing
- |
  shears
- |
  sheath
- |
  sheathe
- |
  sheathing
- |
  sheave
- |
  sheaves
- |
  Sheba
- |
  shebang
- |
  Shebat
- |
  shedder
- |
  shedding
- |
  sheen
- |
  sheeny
- |
  sheep
- |
  sheepcote
- |
  sheepdog
- |
  sheepfold
- |
  sheepish
- |
  sheepishly
- |
  sheepishness
- |
  sheepskin
- |
  sheer
- |
  sheerness
- |
  sheet
- |
  sheeting
- |
  Sheetrock
- |
  sheets
- |
  Sheffield
- |
  sheik
- |
  sheikdom
- |
  sheikh
- |
  sheikhdom
- |
  Sheila
- |
  shekel
- |
  shekels
- |
  Shelby
- |
  Sheldon
- |
  shelf
- |
  Shelia
- |
  shell
- |
  shellac
- |
  shellack
- |
  shellacking
- |
  shelled
- |
  sheller
- |
  Shelley
- |
  shellfire
- |
  shellfish
- |
  shellfishing
- |
  shelling
- |
  shellshocked
- |
  shelly
- |
  shelter
- |
  sheltered
- |
  shelve
- |
  shelves
- |
  shelving
- |
  Shenandoah
- |
  shenanigan
- |
  shenanigans
- |
  Shenyang
- |
  Shepard
- |
  shepherd
- |
  shepherdess
- |
  sheqalim
- |
  sheqel
- |
  sherbert
- |
  sherbet
- |
  Sherbrooke
- |
  sherd
- |
  Sheridan
- |
  sheriff
- |
  Sherman
- |
  Sherpa
- |
  Sherri
- |
  Sherrie
- |
  Sherrill
- |
  Sherry
- |
  sherry
- |
  Sherwin
- |
  Sherwood
- |
  Sheryl
- |
  Shetland
- |
  Shevardnadze
- |
  Shevat
- |
  shiatsu
- |
  shiatzu
- |
  shibboleth
- |
  shied
- |
  shield
- |
  shielder
- |
  shier
- |
  shiest
- |
  shift
- |
  shifter
- |
  shiftily
- |
  shiftiness
- |
  shifting
- |
  shiftless
- |
  shifty
- |
  Shiism
- |
  Shiite
- |
  Shijiazhuang
- |
  Shikoku
- |
  shiksa
- |
  shill
- |
  shillalah
- |
  shillelagh
- |
  shilling
- |
  shimmer
- |
  shimmeringly
- |
  shimmery
- |
  shimmy
- |
  shinbone
- |
  shindig
- |
  shindy
- |
  shine
- |
  shiner
- |
  shingle
- |
  shingler
- |
  shingles
- |
  shingly
- |
  shinguard
- |
  shininess
- |
  shining
- |
  shinny
- |
  shinsplints
- |
  Shinto
- |
  Shintoism
- |
  Shintoist
- |
  shiny
- |
  shipboard
- |
  shipbuilder
- |
  shipbuilding
- |
  shipfitter
- |
  shipload
- |
  shipmaster
- |
  shipmate
- |
  shipment
- |
  shipper
- |
  shipping
- |
  shipshape
- |
  shipworm
- |
  shipwreck
- |
  shipwright
- |
  shipyard
- |
  Shiraz
- |
  shire
- |
  Shires
- |
  shirk
- |
  shirker
- |
  Shirley
- |
  shirr
- |
  shirring
- |
  shirt
- |
  shirtfront
- |
  shirting
- |
  shirtless
- |
  shirtsleeves
- |
  shirttail
- |
  shirtwaist
- |
  shitty
- |
  Shiva
- |
  shiva
- |
  shivah
- |
  shivaree
- |
  shiver
- |
  shiverer
- |
  shivery
- |
  shlemiel
- |
  shlep
- |
  shlepp
- |
  shlock
- |
  shmaltz
- |
  shmear
- |
  shmeer
- |
  shmooze
- |
  shmuck
- |
  shnook
- |
  shnorrer
- |
  Shoah
- |
  shoal
- |
  shoals
- |
  shoat
- |
  shock
- |
  shockability
- |
  shockable
- |
  shocked
- |
  shocker
- |
  shocking
- |
  shockingly
- |
  shockproof
- |
  shockwave
- |
  shodden
- |
  shoddily
- |
  shoddiness
- |
  shoddy
- |
  shoehorn
- |
  shoelace
- |
  shoemaker
- |
  shoemaking
- |
  shoeshine
- |
  shoestring
- |
  shoetree
- |
  shofar
- |
  shofroth
- |
  shogun
- |
  shogunate
- |
  shone
- |
  shook
- |
  shoot
- |
  shooter
- |
  shooting
- |
  shootout
- |
  shopkeeper
- |
  shoplift
- |
  shoplifter
- |
  shoplifting
- |
  shoppe
- |
  shopper
- |
  shopping
- |
  shoptalk
- |
  shopworn
- |
  shore
- |
  shorebird
- |
  shoreless
- |
  shoreline
- |
  shoring
- |
  shorn
- |
  short
- |
  shortage
- |
  shortbread
- |
  shortcake
- |
  shortchange
- |
  shortcoming
- |
  shortcut
- |
  shorten
- |
  shortener
- |
  shortening
- |
  shortfall
- |
  shorthand
- |
  shorthanded
- |
  Shorthorn
- |
  shorthorn
- |
  shortie
- |
  shortish
- |
  shortlist
- |
  shortly
- |
  shortness
- |
  shorts
- |
  shortsighted
- |
  shortstop
- |
  shortwave
- |
  shorty
- |
  Shoshone
- |
  Shoshonean
- |
  Shoshoni
- |
  shotgun
- |
  should
- |
  shoulder
- |
  shoulders
- |
  shout
- |
  shouter
- |
  shove
- |
  shovel
- |
  shovelful
- |
  shover
- |
  Showa
- |
  showbiz
- |
  showboat
- |
  showcase
- |
  showdown
- |
  shower
- |
  showery
- |
  showgirl
- |
  showily
- |
  showiness
- |
  showing
- |
  showman
- |
  showmanship
- |
  shown
- |
  showoff
- |
  showpiece
- |
  showplace
- |
  showroom
- |
  showstopper
- |
  showy
- |
  shrank
- |
  shrapnel
- |
  shred
- |
  shreddable
- |
  shredder
- |
  Shreveport
- |
  shrew
- |
  shrewd
- |
  shrewdly
- |
  shrewdness
- |
  shrewish
- |
  shrewishly
- |
  shrewishness
- |
  Shrewsbury
- |
  shriek
- |
  shrift
- |
  shrike
- |
  shrill
- |
  shrillness
- |
  shrilly
- |
  shrimp
- |
  shrimper
- |
  shrine
- |
  shrink
- |
  shrinkable
- |
  shrinkage
- |
  shrinker
- |
  shrive
- |
  shrivel
- |
  shriveled
- |
  shrivelled
- |
  shriven
- |
  Shropshire
- |
  shroud
- |
  shrouded
- |
  shrove
- |
  shrub
- |
  shrubbery
- |
  shrubbiness
- |
  shrubby
- |
  shrug
- |
  shrunk
- |
  shrunken
- |
  shtick
- |
  shuck
- |
  shucker
- |
  shucks
- |
  shudder
- |
  shudderingly
- |
  shuffle
- |
  shuffleboard
- |
  shuffler
- |
  shunt
- |
  shush
- |
  shutdown
- |
  shuteye
- |
  shutout
- |
  shutter
- |
  shutterbug
- |
  shuttle
- |
  shuttlecock
- |
  shyer
- |
  Shylock
- |
  shylock
- |
  shyly
- |
  shyness
- |
  shyster
- |
  Siamese
- |
  Sibelius
- |
  Siberia
- |
  Siberian
- |
  sibilance
- |
  sibilancy
- |
  sibilant
- |
  sibilantly
- |
  sibilate
- |
  sibilation
- |
  sibling
- |
  Sibyl
- |
  sibyl
- |
  sibylline
- |
  Sichuan
- |
  Sicilian
- |
  Sicily
- |
  sickbay
- |
  sickbed
- |
  sicken
- |
  sickening
- |
  sickeningly
- |
  sickie
- |
  sickish
- |
  sickle
- |
  sickliness
- |
  sickly
- |
  sickness
- |
  sicko
- |
  sickout
- |
  sickroom
- |
  Siddhartha
- |
  sidearm
- |
  sidebar
- |
  sideboard
- |
  sideburns
- |
  sidecar
- |
  sidekick
- |
  sidelight
- |
  sideline
- |
  sidelong
- |
  sideman
- |
  sidepiece
- |
  sidereal
- |
  sidesaddle
- |
  sideshow
- |
  sideslip
- |
  sidestep
- |
  sidestroke
- |
  sideswipe
- |
  sidetrack
- |
  sidewalk
- |
  sidewall
- |
  sideways
- |
  sidewinder
- |
  sidewise
- |
  siding
- |
  sidle
- |
  Sidney
- |
  Sidon
- |
  siege
- |
  Siegfried
- |
  Siemens
- |
  siemens
- |
  Siena
- |
  Sienese
- |
  sienna
- |
  sierra
- |
  sierran
- |
  siesta
- |
  sieve
- |
  sifter
- |
  sigher
- |
  sight
- |
  sighted
- |
  sighting
- |
  sightless
- |
  sightlessly
- |
  sightliness
- |
  sightly
- |
  sightread
- |
  sightseeing
- |
  sightseer
- |
  sigil
- |
  sigma
- |
  Sigmund
- |
  signage
- |
  signal
- |
  signaler
- |
  signalize
- |
  signaller
- |
  signally
- |
  signalman
- |
  signatory
- |
  signature
- |
  signboard
- |
  signer
- |
  signet
- |
  significance
- |
  significant
- |
  signifier
- |
  signify
- |
  signing
- |
  signor
- |
  signora
- |
  signore
- |
  signori
- |
  signorina
- |
  signorine
- |
  signpost
- |
  Sigrid
- |
  Sikhism
- |
  Sikkim
- |
  Sikorsky
- |
  silage
- |
  Silas
- |
  silence
- |
  silencer
- |
  sileni
- |
  silent
- |
  silently
- |
  Silenus
- |
  silenus
- |
  Silesia
- |
  Silesian
- |
  silhouette
- |
  silica
- |
  silicate
- |
  siliceous
- |
  silicious
- |
  silicon
- |
  silicone
- |
  silicosis
- |
  silken
- |
  silkily
- |
  silkiness
- |
  silkscreen
- |
  silkworm
- |
  silky
- |
  silliness
- |
  silly
- |
  siltation
- |
  silty
- |
  Silurian
- |
  silvan
- |
  silver
- |
  silverer
- |
  silverfish
- |
  silveriness
- |
  silversmith
- |
  silverware
- |
  silvery
- |
  Silvester
- |
  Silvia
- |
  silviculture
- |
  Simbirsk
- |
  Simeon
- |
  Simferopol
- |
  simian
- |
  similar
- |
  similarity
- |
  similarly
- |
  simile
- |
  similitude
- |
  simmer
- |
  Simon
- |
  simoniac
- |
  simoniacal
- |
  simonize
- |
  simony
- |
  simpatico
- |
  simper
- |
  simperer
- |
  simperingly
- |
  simple
- |
  simpleness
- |
  simpleton
- |
  simplicity
- |
  simplified
- |
  simplifier
- |
  simplify
- |
  simplism
- |
  simplistic
- |
  simply
- |
  simulacra
- |
  simulacrum
- |
  simulate
- |
  simulated
- |
  simulation
- |
  simulative
- |
  simulator
- |
  simulcast
- |
  simultaneity
- |
  simultaneous
- |
  Sinai
- |
  Sinaloa
- |
  Sinatra
- |
  since
- |
  sincere
- |
  sincerely
- |
  sincereness
- |
  sincerity
- |
  Sinclair
- |
  Sindbad
- |
  sinecure
- |
  sinecurism
- |
  sinecurist
- |
  sinew
- |
  sinewed
- |
  sinews
- |
  sinewy
- |
  sinfonia
- |
  sinfonietta
- |
  sinful
- |
  sinfully
- |
  sinfulness
- |
  singable
- |
  Singapore
- |
  Singaporean
- |
  singe
- |
  Singer
- |
  singer
- |
  Singhalese
- |
  singing
- |
  single
- |
  singleness
- |
  singles
- |
  singleton
- |
  singletree
- |
  singly
- |
  singsong
- |
  singspiel
- |
  singspiele
- |
  singular
- |
  singularity
- |
  singularly
- |
  singularness
- |
  Sinhalese
- |
  sinister
- |
  sinisterly
- |
  sinisterness
- |
  sinistral
- |
  sinistrality
- |
  sinistrally
- |
  sinkable
- |
  sinker
- |
  sinkhole
- |
  sinking
- |
  sinless
- |
  sinner
- |
  Sinologist
- |
  Sinology
- |
  sinter
- |
  sinuosity
- |
  sinuous
- |
  sinuously
- |
  sinuousness
- |
  sinus
- |
  sinusitis
- |
  Siouan
- |
  Sioux
- |
  siphon
- |
  sipper
- |
  Sirach
- |
  siree
- |
  Siren
- |
  siren
- |
  Sirius
- |
  sirloin
- |
  sirocco
- |
  sirree
- |
  sirup
- |
  sisal
- |
  sissified
- |
  sissy
- |
  sissyish
- |
  Sister
- |
  sister
- |
  sisterhood
- |
  sisterliness
- |
  sisterly
- |
  Sisyphean
- |
  Sisyphus
- |
  sitar
- |
  sitarist
- |
  sitcom
- |
  siting
- |
  sitter
- |
  sitting
- |
  situate
- |
  situated
- |
  situation
- |
  situational
- |
  situationism
- |
  situationist
- |
  situp
- |
  situs
- |
  Sivan
- |
  sixpence
- |
  sixteen
- |
  sixteenth
- |
  sixth
- |
  sixtieth
- |
  sixty
- |
  sizable
- |
  sizableness
- |
  sizably
- |
  sizeable
- |
  sized
- |
  sizing
- |
  sizzle
- |
  sizzlingly
- |
  Sjaelland
- |
  Skagerak
- |
  Skagerrak
- |
  Skagway
- |
  skald
- |
  skaldic
- |
  skate
- |
  skateboard
- |
  skateboarder
- |
  skater
- |
  skating
- |
  skedaddle
- |
  skeet
- |
  skein
- |
  skeletal
- |
  skeleton
- |
  skeptic
- |
  skeptical
- |
  skeptically
- |
  skepticism
- |
  sketch
- |
  sketcher
- |
  sketchily
- |
  sketchiness
- |
  sketchy
- |
  skewbald
- |
  skewed
- |
  skewer
- |
  skewness
- |
  skiable
- |
  skids
- |
  skier
- |
  skies
- |
  skiff
- |
  skiing
- |
  skilful
- |
  skilfully
- |
  skill
- |
  skilled
- |
  skillet
- |
  skillful
- |
  skillfully
- |
  skillfulness
- |
  skimmer
- |
  skimp
- |
  skimpily
- |
  skimpiness
- |
  skimpy
- |
  skincare
- |
  skinflick
- |
  skinflint
- |
  skinhead
- |
  skinless
- |
  skinned
- |
  Skinner
- |
  skinniness
- |
  skinny
- |
  skintight
- |
  skipjack
- |
  skipper
- |
  skipping
- |
  skirmish
- |
  skirmishing
- |
  skirt
- |
  skitter
- |
  skittish
- |
  skittishly
- |
  skittishness
- |
  skivvies
- |
  skivvy
- |
  skiwear
- |
  skoal
- |
  Skopje
- |
  Skoplje
- |
  skosh
- |
  skulduggery
- |
  skulk
- |
  skulker
- |
  skull
- |
  skullcap
- |
  skullduggery
- |
  skunk
- |
  skycap
- |
  skydive
- |
  skydiver
- |
  skydiving
- |
  skyhook
- |
  skyjack
- |
  skyjacker
- |
  skyjacking
- |
  skylark
- |
  skylight
- |
  skylighted
- |
  skyline
- |
  skyrocket
- |
  skyscraper
- |
  skywalk
- |
  skyward
- |
  skywards
- |
  skywriter
- |
  skywriting
- |
  slack
- |
  slacken
- |
  slackening
- |
  slacker
- |
  slackly
- |
  slackness
- |
  slacks
- |
  slagging
- |
  slaggy
- |
  slain
- |
  slake
- |
  slalom
- |
  slammer
- |
  slander
- |
  slanderer
- |
  slanderous
- |
  slanderously
- |
  slang
- |
  slanginess
- |
  slangy
- |
  slant
- |
  slanted
- |
  slantingly
- |
  slantwise
- |
  slapdash
- |
  slaphappy
- |
  slapstick
- |
  slash
- |
  slasher
- |
  slate
- |
  slather
- |
  slattern
- |
  slatternly
- |
  slaty
- |
  slaughter
- |
  slaughterer
- |
  slave
- |
  slaver
- |
  slavery
- |
  Slavic
- |
  slavish
- |
  slavishly
- |
  slavishness
- |
  Slavonia
- |
  Slavonian
- |
  Slavonic
- |
  slayer
- |
  slaying
- |
  sleaze
- |
  sleazily
- |
  sleaziness
- |
  sleazy
- |
  sledder
- |
  sledge
- |
  sledgehammer
- |
  sleek
- |
  sleekly
- |
  sleekness
- |
  sleep
- |
  sleeper
- |
  sleepily
- |
  sleepiness
- |
  sleepless
- |
  sleeplessly
- |
  sleepwalk
- |
  sleepwalker
- |
  sleepwalking
- |
  sleepwear
- |
  sleepy
- |
  sleepyhead
- |
  sleet
- |
  sleety
- |
  sleeve
- |
  sleeved
- |
  sleeveless
- |
  sleigh
- |
  sleight
- |
  slender
- |
  slenderize
- |
  slenderly
- |
  slenderness
- |
  slept
- |
  sleuth
- |
  sleuthhound
- |
  sleuthing
- |
  slice
- |
  sliceable
- |
  slicer
- |
  slick
- |
  slicker
- |
  slickly
- |
  slickness
- |
  slide
- |
  slider
- |
  slier
- |
  sliest
- |
  slight
- |
  slighting
- |
  slightly
- |
  slightness
- |
  slily
- |
  slime
- |
  sliminess
- |
  slimly
- |
  slimmer
- |
  slimming
- |
  slimmish
- |
  slimness
- |
  slimy
- |
  sling
- |
  slinger
- |
  slingshot
- |
  slink
- |
  slinkily
- |
  slinkiness
- |
  slinky
- |
  slipcase
- |
  slipcover
- |
  slipknot
- |
  slippage
- |
  slipper
- |
  slipperiness
- |
  slippery
- |
  slipshod
- |
  slipstream
- |
  slipup
- |
  slither
- |
  slithery
- |
  sliver
- |
  slobber
- |
  slobberer
- |
  slogan
- |
  sloop
- |
  slope
- |
  sloping
- |
  sloppily
- |
  sloppiness
- |
  sloppy
- |
  slops
- |
  slosh
- |
  sloshed
- |
  sloshy
- |
  sloth
- |
  slothful
- |
  slothfully
- |
  slothfulness
- |
  slouch
- |
  slouched
- |
  sloucher
- |
  slouchy
- |
  slough
- |
  sloughy
- |
  Slovak
- |
  Slovakia
- |
  Slovakian
- |
  sloven
- |
  Slovene
- |
  Slovenia
- |
  Slovenian
- |
  slovenliness
- |
  slovenly
- |
  slowdown
- |
  slowly
- |
  slowness
- |
  slowpoke
- |
  sludge
- |
  sludgy
- |
  sluff
- |
  sluggard
- |
  sluggardly
- |
  slugger
- |
  sluggish
- |
  sluggishly
- |
  sluggishness
- |
  sluice
- |
  sluiceway
- |
  slumber
- |
  slumberer
- |
  slumberous
- |
  slumbrous
- |
  slumlord
- |
  slummy
- |
  slump
- |
  slung
- |
  slunk
- |
  slurp
- |
  slurred
- |
  slurry
- |
  slush
- |
  slushily
- |
  slushiness
- |
  slushy
- |
  sluttish
- |
  slyly
- |
  slyness
- |
  smack
- |
  smacker
- |
  small
- |
  smallish
- |
  smallness
- |
  smallpox
- |
  smalltime
- |
  smalltimer
- |
  smarmily
- |
  smarminess
- |
  smarmy
- |
  smart
- |
  smarten
- |
  smartly
- |
  smartness
- |
  smarts
- |
  smash
- |
  smashed
- |
  smasher
- |
  smashing
- |
  smashup
- |
  smatter
- |
  smattering
- |
  smear
- |
  smeared
- |
  smeary
- |
  smegma
- |
  smell
- |
  smelliness
- |
  smelly
- |
  smelt
- |
  smelter
- |
  smeltery
- |
  smelting
- |
  Smetana
- |
  smidge
- |
  smidgen
- |
  smidgeon
- |
  smidgin
- |
  smilax
- |
  smile
- |
  smiley
- |
  smilingly
- |
  smirch
- |
  smirk
- |
  smirker
- |
  smirkily
- |
  smirkingly
- |
  smirky
- |
  smite
- |
  smiter
- |
  Smith
- |
  smith
- |
  smithereens
- |
  Smithson
- |
  smithy
- |
  smitten
- |
  smock
- |
  smocking
- |
  smoggy
- |
  smoke
- |
  smokehouse
- |
  smokeless
- |
  smoker
- |
  smokescreen
- |
  smokestack
- |
  smokiness
- |
  smoking
- |
  smoky
- |
  smolder
- |
  smoldering
- |
  smolderingly
- |
  Smolensk
- |
  Smollett
- |
  smooch
- |
  smooth
- |
  smoothbore
- |
  smoother
- |
  smoothie
- |
  smoothly
- |
  smoothness
- |
  smorgasbord
- |
  smote
- |
  smother
- |
  smothered
- |
  smoulder
- |
  smudge
- |
  smudgy
- |
  smuggle
- |
  smuggler
- |
  smuggling
- |
  smugly
- |
  smugness
- |
  smutch
- |
  Smuts
- |
  smuttiness
- |
  smutty
- |
  Smyrna
- |
  snack
- |
  snaffle
- |
  snafu
- |
  snail
- |
  Snake
- |
  snake
- |
  snakebite
- |
  snakelike
- |
  snakily
- |
  snaky
- |
  snapdragon
- |
  snapper
- |
  snappily
- |
  snappish
- |
  snappy
- |
  snapshot
- |
  snare
- |
  snarl
- |
  snarler
- |
  snarlingly
- |
  snarly
- |
  snatch
- |
  snatcher
- |
  snazzily
- |
  snazziness
- |
  snazzy
- |
  sneak
- |
  sneaker
- |
  sneakily
- |
  sneakiness
- |
  sneaking
- |
  sneakingly
- |
  sneaky
- |
  sneer
- |
  sneering
- |
  sneeringly
- |
  sneeze
- |
  snicker
- |
  snickeringly
- |
  snide
- |
  snidely
- |
  snideness
- |
  snidey
- |
  sniff
- |
  sniffer
- |
  sniffle
- |
  sniffles
- |
  snifter
- |
  snigger
- |
  sniggerer
- |
  sniggeringly
- |
  snipe
- |
  sniper
- |
  snippet
- |
  snippiness
- |
  snippy
- |
  snips
- |
  snitch
- |
  snivel
- |
  sniveler
- |
  sniveling
- |
  snivelingly
- |
  snobbery
- |
  snobbish
- |
  snobbishly
- |
  snobbishness
- |
  snobby
- |
  snood
- |
  snooker
- |
  snoop
- |
  snooper
- |
  snoopily
- |
  snoopiness
- |
  snoopy
- |
  snoot
- |
  snootful
- |
  snootily
- |
  snootiness
- |
  snooty
- |
  snooze
- |
  snoozer
- |
  snore
- |
  snorer
- |
  snorkel
- |
  snorkeler
- |
  snorkeling
- |
  snort
- |
  snorter
- |
  snottily
- |
  snottiness
- |
  snotty
- |
  snout
- |
  snowball
- |
  snowbank
- |
  Snowbelt
- |
  snowbelt
- |
  snowblower
- |
  snowboard
- |
  snowboarder
- |
  snowboarding
- |
  snowbound
- |
  Snowdon
- |
  Snowdonia
- |
  snowdrift
- |
  snowdrop
- |
  snowfall
- |
  snowfield
- |
  snowflake
- |
  snowman
- |
  snowmobile
- |
  snowmobiler
- |
  snowmobiling
- |
  snowplow
- |
  snowshoe
- |
  snowstorm
- |
  snowsuit
- |
  snowy
- |
  snuck
- |
  snuff
- |
  snuffbox
- |
  snuffer
- |
  snuffle
- |
  snuffler
- |
  snuffling
- |
  snuffly
- |
  snuggle
- |
  snugly
- |
  snugness
- |
  soaked
- |
  soaker
- |
  soaking
- |
  soapbox
- |
  soapily
- |
  soapiness
- |
  soapstone
- |
  soapsuds
- |
  soapy
- |
  soaring
- |
  Soave
- |
  sobbing
- |
  sobbingly
- |
  sober
- |
  sobering
- |
  soberly
- |
  soberness
- |
  sobriety
- |
  sobriquet
- |
  soccer
- |
  sociability
- |
  sociable
- |
  sociableness
- |
  sociably
- |
  social
- |
  socialise
- |
  socialism
- |
  socialist
- |
  socialistic
- |
  socialite
- |
  sociality
- |
  socialize
- |
  socializer
- |
  socializing
- |
  socially
- |
  societal
- |
  Society
- |
  society
- |
  sociobiology
- |
  sociologic
- |
  sociological
- |
  sociologist
- |
  sociology
- |
  sociometric
- |
  sociometrist
- |
  sociometry
- |
  sociopath
- |
  sociopathic
- |
  sociopathy
- |
  socket
- |
  Socotra
- |
  Socrates
- |
  Socratic
- |
  sodality
- |
  sodden
- |
  soddenly
- |
  soddenness
- |
  sodium
- |
  Sodom
- |
  sodomite
- |
  sodomize
- |
  sodomy
- |
  soever
- |
  sofabed
- |
  soffit
- |
  Sofia
- |
  softball
- |
  softbound
- |
  soften
- |
  softener
- |
  softhearted
- |
  softie
- |
  softly
- |
  softness
- |
  software
- |
  softwood
- |
  softy
- |
  soggily
- |
  sogginess
- |
  soggy
- |
  soigne
- |
  soignee
- |
  soiled
- |
  soiree
- |
  sojourn
- |
  sojourner
- |
  solace
- |
  solacer
- |
  solar
- |
  solaria
- |
  solarium
- |
  solder
- |
  solderer
- |
  soldier
- |
  soldiering
- |
  soldierly
- |
  soldiery
- |
  solecism
- |
  solecistic
- |
  solely
- |
  solemn
- |
  solemness
- |
  solemnities
- |
  solemnity
- |
  solemnize
- |
  solemnly
- |
  solemnness
- |
  solenoid
- |
  soles
- |
  solicit
- |
  solicitation
- |
  soliciting
- |
  solicitor
- |
  solicitous
- |
  solicitously
- |
  solicitude
- |
  solid
- |
  Solidarity
- |
  solidarity
- |
  solidi
- |
  solidify
- |
  solidity
- |
  solidly
- |
  solidness
- |
  solids
- |
  solidus
- |
  Solihull
- |
  soliloquist
- |
  soliloquize
- |
  soliloquy
- |
  solipsism
- |
  solipsist
- |
  solipsistic
- |
  solitaire
- |
  solitarily
- |
  solitariness
- |
  solitary
- |
  solitude
- |
  solmization
- |
  soloist
- |
  Solomon
- |
  Solon
- |
  solon
- |
  Solonian
- |
  Solonic
- |
  solstice
- |
  solstitial
- |
  solubility
- |
  soluble
- |
  solubly
- |
  solute
- |
  solution
- |
  solvable
- |
  solve
- |
  solvency
- |
  solvent
- |
  solver
- |
  Solzhenitsyn
- |
  Somali
- |
  Somalia
- |
  Somalian
- |
  Somaliland
- |
  somatic
- |
  somatically
- |
  somatotype
- |
  somatotyping
- |
  somber
- |
  somberly
- |
  somberness
- |
  sombre
- |
  sombrely
- |
  sombrero
- |
  somebody
- |
  someday
- |
  somehow
- |
  someone
- |
  someplace
- |
  somersault
- |
  Somerset
- |
  somerset
- |
  something
- |
  sometime
- |
  sometimes
- |
  someway
- |
  someways
- |
  somewhat
- |
  somewhere
- |
  Somme
- |
  sommelier
- |
  somnambulant
- |
  somnambulate
- |
  somnambulism
- |
  somnambulist
- |
  somniferous
- |
  somnolence
- |
  somnolency
- |
  somnolent
- |
  somnolently
- |
  sonant
- |
  sonar
- |
  sonata
- |
  sonatina
- |
  Sondheim
- |
  Sondra
- |
  songbird
- |
  songfest
- |
  Songhua
- |
  songster
- |
  songstress
- |
  songwriter
- |
  Sonia
- |
  sonic
- |
  sonically
- |
  sonics
- |
  Sonja
- |
  sonly
- |
  sonnet
- |
  sonny
- |
  sonogram
- |
  Sonora
- |
  Sonoran
- |
  sonority
- |
  sonorous
- |
  sonorously
- |
  sonorousness
- |
  Sonya
- |
  Soochow
- |
  sooner
- |
  sooth
- |
  soothe
- |
  soother
- |
  soothing
- |
  soothingly
- |
  soothsayer
- |
  soothsaying
- |
  sootiness
- |
  sooty
- |
  Sophia
- |
  sophism
- |
  sophist
- |
  sophistic
- |
  sophistical
- |
  sophisticate
- |
  sophistry
- |
  Sophoclean
- |
  Sophocles
- |
  sophomore
- |
  sophomoric
- |
  Sophonias
- |
  soporiferous
- |
  soporific
- |
  soppily
- |
  soppiness
- |
  sopping
- |
  soppy
- |
  sopranino
- |
  soprano
- |
  sorbet
- |
  Sorbian
- |
  sorbitol
- |
  sorcerer
- |
  sorceress
- |
  sorcery
- |
  sordid
- |
  sordidly
- |
  sordidness
- |
  sorehead
- |
  sorely
- |
  soreness
- |
  sorghum
- |
  sororal
- |
  sororicide
- |
  sorority
- |
  sorrel
- |
  sorrily
- |
  sorriness
- |
  sorrow
- |
  sorrowful
- |
  sorrowfully
- |
  sorry
- |
  sorta
- |
  sorter
- |
  sortie
- |
  sortilege
- |
  sostenuto
- |
  soteriology
- |
  sottish
- |
  sottishly
- |
  soubrette
- |
  soubriquet
- |
  souffle
- |
  sough
- |
  sought
- |
  souled
- |
  soulful
- |
  soulfully
- |
  soulfulness
- |
  soulless
- |
  sound
- |
  soundable
- |
  soundboard
- |
  sounder
- |
  sounding
- |
  soundless
- |
  soundlessly
- |
  soundly
- |
  soundness
- |
  soundproof
- |
  soundstage
- |
  soundtrack
- |
  soupcon
- |
  soupy
- |
  sourball
- |
  source
- |
  sourcing
- |
  sourdough
- |
  sourish
- |
  sourly
- |
  sourness
- |
  sourpuss
- |
  soursop
- |
  Sousa
- |
  souse
- |
  soused
- |
  Souter
- |
  South
- |
  south
- |
  Southampton
- |
  southbound
- |
  Southeast
- |
  southeast
- |
  southeaster
- |
  southeastern
- |
  southerly
- |
  southern
- |
  Southerner
- |
  southerner
- |
  southernmost
- |
  Southey
- |
  southpaw
- |
  southward
- |
  southwardly
- |
  southwards
- |
  Southwark
- |
  Southwest
- |
  southwest
- |
  southwester
- |
  southwestern
- |
  souvenir
- |
  sovereign
- |
  sovereignly
- |
  sovereignty
- |
  Soviet
- |
  soviet
- |
  sovietism
- |
  Sovietize
- |
  sovietize
- |
  Soviets
- |
  sower
- |
  Soweto
- |
  soybean
- |
  Soyinka
- |
  soymilk
- |
  space
- |
  spacecraft
- |
  spaced
- |
  spaceflight
- |
  spaceman
- |
  spaceport
- |
  spacer
- |
  spaceship
- |
  spacesuit
- |
  spacewalk
- |
  spacewalker
- |
  spacewoman
- |
  spacey
- |
  spaciness
- |
  spacing
- |
  spacious
- |
  spaciously
- |
  spaciousness
- |
  Spackle
- |
  spacy
- |
  spade
- |
  spadeful
- |
  spader
- |
  spadework
- |
  spadices
- |
  spadix
- |
  spaghetti
- |
  Spain
- |
  spake
- |
  spandex
- |
  spandrel
- |
  spangle
- |
  spangled
- |
  Spanglish
- |
  spangly
- |
  Spaniard
- |
  spaniel
- |
  Spanish
- |
  spank
- |
  spanker
- |
  spanking
- |
  spanner
- |
  spare
- |
  sparely
- |
  spareness
- |
  spareribs
- |
  sparge
- |
  sparger
- |
  sparing
- |
  sparingly
- |
  sparingness
- |
  spark
- |
  sparker
- |
  sparkle
- |
  sparkler
- |
  sparkling
- |
  sparky
- |
  sparrow
- |
  sparse
- |
  sparsely
- |
  sparseness
- |
  sparsity
- |
  Sparta
- |
  Spartacus
- |
  Spartan
- |
  spartan
- |
  spasm
- |
  spasmodic
- |
  spastic
- |
  spastically
- |
  spasticity
- |
  spate
- |
  spathe
- |
  spatial
- |
  spatially
- |
  spatter
- |
  spatula
- |
  spavin
- |
  spavined
- |
  spawn
- |
  spawner
- |
  speak
- |
  speakable
- |
  speakeasy
- |
  speaker
- |
  speaking
- |
  spear
- |
  spearer
- |
  spearfish
- |
  spearfisher
- |
  spearfishing
- |
  spearhead
- |
  spearman
- |
  spearmint
- |
  special
- |
  specialise
- |
  specialised
- |
  specialist
- |
  speciality
- |
  specialize
- |
  specialized
- |
  specially
- |
  specialty
- |
  specie
- |
  species
- |
  speciesism
- |
  speciesist
- |
  specific
- |
  specifically
- |
  specificity
- |
  specifics
- |
  specify
- |
  specimen
- |
  specious
- |
  speciously
- |
  speciousness
- |
  speck
- |
  speckle
- |
  speckled
- |
  specs
- |
  spectacle
- |
  spectacled
- |
  spectacles
- |
  spectacular
- |
  spectator
- |
  specter
- |
  spectra
- |
  spectral
- |
  spectrally
- |
  spectre
- |
  spectrogram
- |
  spectrograph
- |
  spectrometer
- |
  spectrometry
- |
  spectroscope
- |
  spectroscopy
- |
  spectrum
- |
  specula
- |
  specular
- |
  speculate
- |
  speculation
- |
  speculative
- |
  speculator
- |
  speculum
- |
  speech
- |
  speechless
- |
  speechlessly
- |
  speed
- |
  speedboat
- |
  speeder
- |
  speedily
- |
  speediness
- |
  speeding
- |
  speedometer
- |
  speedster
- |
  speedup
- |
  speedway
- |
  speedwell
- |
  speedy
- |
  speleologist
- |
  speleology
- |
  spell
- |
  spellbind
- |
  spellbinder
- |
  spellbinding
- |
  spellbound
- |
  spelldown
- |
  speller
- |
  spelling
- |
  spelt
- |
  spelunker
- |
  spelunking
- |
  Spencer
- |
  spend
- |
  spendable
- |
  spender
- |
  spending
- |
  spendthrift
- |
  Spenser
- |
  Spenserian
- |
  spent
- |
  sperm
- |
  spermaceti
- |
  spermatic
- |
  spermatozoa
- |
  spermatozoon
- |
  spermicidal
- |
  spermicide
- |
  spewer
- |
  sphagnum
- |
  sphere
- |
  spherical
- |
  spherically
- |
  spheroid
- |
  spheroidal
- |
  sphincter
- |
  sphincteral
- |
  sphincteric
- |
  sphinges
- |
  Sphinx
- |
  sphinx
- |
  sphinxlike
- |
  Spica
- |
  spice
- |
  spiced
- |
  spiciness
- |
  spicule
- |
  spicy
- |
  spider
- |
  spiderweb
- |
  spidery
- |
  spiel
- |
  Spielberg
- |
  spiffily
- |
  spiffy
- |
  spigot
- |
  spike
- |
  spiked
- |
  spikelet
- |
  spikenard
- |
  spiky
- |
  spill
- |
  spillable
- |
  spillage
- |
  spillway
- |
  spilt
- |
  spinach
- |
  spinal
- |
  spinally
- |
  spindle
- |
  spindling
- |
  spindly
- |
  spindrift
- |
  spine
- |
  spinel
- |
  spineless
- |
  spinet
- |
  spinnaker
- |
  spinner
- |
  spinneret
- |
  spinning
- |
  spinoff
- |
  Spinoza
- |
  spinster
- |
  spinsterhood
- |
  spinsterish
- |
  spiny
- |
  spiracle
- |
  spiraea
- |
  spiral
- |
  spirally
- |
  spirant
- |
  spire
- |
  spirea
- |
  Spirit
- |
  spirit
- |
  spirited
- |
  spiritedly
- |
  spiritless
- |
  spirits
- |
  spiritual
- |
  spiritualism
- |
  spiritualist
- |
  spirituality
- |
  spiritualize
- |
  spiritually
- |
  spirituous
- |
  spirochaete
- |
  spirochete
- |
  spirt
- |
  spiry
- |
  spitball
- |
  spite
- |
  spiteful
- |
  spitefully
- |
  spitefulness
- |
  spitfire
- |
  spittle
- |
  spittlebug
- |
  spittoon
- |
  splash
- |
  splashdown
- |
  splasher
- |
  splashily
- |
  splashiness
- |
  splashy
- |
  splat
- |
  splatter
- |
  splay
- |
  splayed
- |
  splayfeet
- |
  splayfoot
- |
  splayfooted
- |
  spleen
- |
  spleenful
- |
  splendent
- |
  splendid
- |
  splendidly
- |
  splendor
- |
  splendorous
- |
  splendour
- |
  splendrous
- |
  splenetic
- |
  splenic
- |
  splice
- |
  splicer
- |
  spline
- |
  splined
- |
  splint
- |
  splinter
- |
  splintery
- |
  Split
- |
  split
- |
  splitter
- |
  splitting
- |
  splotch
- |
  splotchy
- |
  splurge
- |
  splutter
- |
  Spock
- |
  spoil
- |
  spoilage
- |
  spoiled
- |
  spoiler
- |
  spoils
- |
  spoilsport
- |
  spoilt
- |
  Spokane
- |
  spoke
- |
  spoken
- |
  spokesman
- |
  spokespeople
- |
  spokesperson
- |
  spokeswoman
- |
  spoliation
- |
  spoliator
- |
  spondaic
- |
  spondee
- |
  sponge
- |
  spongecake
- |
  sponger
- |
  spongiform
- |
  sponginess
- |
  spongy
- |
  sponsor
- |
  sponsored
- |
  sponsorship
- |
  spontaneity
- |
  spontaneous
- |
  spoof
- |
  spook
- |
  spooked
- |
  spookily
- |
  spookiness
- |
  spooky
- |
  spool
- |
  spooler
- |
  spoon
- |
  spoonbill
- |
  spoonerism
- |
  spoonfed
- |
  spoonfeed
- |
  spoonful
- |
  spoor
- |
  spoorer
- |
  Sporades
- |
  sporadic
- |
  sporadically
- |
  spore
- |
  sporran
- |
  sport
- |
  sportily
- |
  sportiness
- |
  sporting
- |
  sportingly
- |
  sportive
- |
  sportively
- |
  sportiveness
- |
  sports
- |
  sportscast
- |
  sportscaster
- |
  sportsman
- |
  sportswear
- |
  sportswoman
- |
  sportswriter
- |
  sporty
- |
  spotless
- |
  spotlessly
- |
  spotlessness
- |
  spotlight
- |
  spotted
- |
  spotter
- |
  spottily
- |
  spottiness
- |
  spotty
- |
  spousal
- |
  spousals
- |
  spouse
- |
  spout
- |
  spouter
- |
  sprain
- |
  sprang
- |
  sprat
- |
  sprawl
- |
  sprawled
- |
  spray
- |
  sprayer
- |
  spread
- |
  spreadable
- |
  spreader
- |
  spreadsheet
- |
  Sprechgesang
- |
  sprechgesang
- |
  spree
- |
  sprier
- |
  spriest
- |
  sprig
- |
  sprightly
- |
  spring
- |
  springboard
- |
  springe
- |
  Springfield
- |
  springily
- |
  springiness
- |
  springlike
- |
  Springsteen
- |
  springtime
- |
  springy
- |
  sprinkle
- |
  sprinkler
- |
  sprinkling
- |
  sprint
- |
  sprinter
- |
  sprite
- |
  spritz
- |
  spritzer
- |
  sprocket
- |
  sprout
- |
  spruce
- |
  sprucely
- |
  spruceness
- |
  sprung
- |
  spryly
- |
  spryness
- |
  spume
- |
  spumone
- |
  spumoni
- |
  spumous
- |
  spumy
- |
  spunk
- |
  spunky
- |
  spurge
- |
  spurious
- |
  spuriously
- |
  spuriousness
- |
  spurn
- |
  spurner
- |
  spurred
- |
  spurt
- |
  sputa
- |
  Sputnik
- |
  sputnik
- |
  sputter
- |
  sputterer
- |
  sputum
- |
  spyglass
- |
  spying
- |
  squab
- |
  squabble
- |
  squabbler
- |
  squad
- |
  squadron
- |
  squalid
- |
  squalidly
- |
  squalidness
- |
  squall
- |
  squally
- |
  squalor
- |
  squamose
- |
  squamous
- |
  squander
- |
  squanderer
- |
  Squanto
- |
  square
- |
  squarely
- |
  squareness
- |
  squarish
- |
  squash
- |
  squashiness
- |
  squashy
- |
  squat
- |
  squatness
- |
  squatter
- |
  squaw
- |
  squawk
- |
  squeak
- |
  squeaker
- |
  squeakily
- |
  squeakiness
- |
  squeaky
- |
  squeal
- |
  squealer
- |
  squeamish
- |
  squeamishly
- |
  squeegee
- |
  squeezable
- |
  squeeze
- |
  squeezer
- |
  squelch
- |
  squelcher
- |
  squelchy
- |
  squib
- |
  squibber
- |
  squid
- |
  squiggle
- |
  squiggly
- |
  squint
- |
  squinty
- |
  squire
- |
  squiredom
- |
  squireship
- |
  squirm
- |
  squirmer
- |
  squirmy
- |
  squirrel
- |
  squirt
- |
  squish
- |
  squishy
- |
  Srinagar
- |
  stabbing
- |
  stabile
- |
  stabilise
- |
  stability
- |
  stabilize
- |
  stabilizer
- |
  stable
- |
  stableman
- |
  stably
- |
  staccato
- |
  Stacey
- |
  stack
- |
  stacker
- |
  stacks
- |
  stackup
- |
  Stacy
- |
  stadia
- |
  stadium
- |
  Stael
- |
  staff
- |
  staffed
- |
  staffer
- |
  staffing
- |
  Stafford
- |
  stage
- |
  stageable
- |
  stagecoach
- |
  stagecraft
- |
  stagefright
- |
  stagehand
- |
  stagestruck
- |
  stagey
- |
  stagflation
- |
  stagger
- |
  staggered
- |
  staggerer
- |
  staggering
- |
  staggeringly
- |
  staggers
- |
  stagily
- |
  staginess
- |
  staging
- |
  stagnancy
- |
  stagnant
- |
  stagnantly
- |
  stagnate
- |
  stagnation
- |
  stagy
- |
  staid
- |
  staidly
- |
  staidness
- |
  stain
- |
  stained
- |
  stainless
- |
  stair
- |
  staircase
- |
  stairs
- |
  stairway
- |
  stairwell
- |
  stake
- |
  stakeout
- |
  stakes
- |
  stalactite
- |
  stalactitic
- |
  Stalag
- |
  stalagmite
- |
  stalagmitic
- |
  stale
- |
  stalely
- |
  stalemate
- |
  stalemated
- |
  staleness
- |
  Stalin
- |
  Stalingrad
- |
  Stalinism
- |
  Stalinist
- |
  stalk
- |
  stalked
- |
  stalker
- |
  stalking
- |
  stall
- |
  stallion
- |
  stalwart
- |
  stalwartly
- |
  stalwartness
- |
  stamen
- |
  Stamford
- |
  stamina
- |
  staminate
- |
  stammer
- |
  stammerer
- |
  stammering
- |
  stammeringly
- |
  stamp
- |
  stampede
- |
  stamper
- |
  stance
- |
  stanch
- |
  stanchion
- |
  stanchioned
- |
  stand
- |
  standalone
- |
  standard
- |
  standardise
- |
  standardize
- |
  standby
- |
  standbys
- |
  standee
- |
  stander
- |
  standing
- |
  Standish
- |
  standoff
- |
  standoffish
- |
  standout
- |
  standpipe
- |
  standpoint
- |
  stands
- |
  standstill
- |
  standup
- |
  Stanford
- |
  Stanislavsky
- |
  stank
- |
  Stanley
- |
  Stanton
- |
  stanza
- |
  stanzaed
- |
  stanzaic
- |
  stapedes
- |
  stapes
- |
  staph
- |
  staple
- |
  stapler
- |
  starboard
- |
  starch
- |
  starchily
- |
  starchiness
- |
  starchy
- |
  stardom
- |
  stardust
- |
  stare
- |
  starer
- |
  starfish
- |
  stargaze
- |
  stargazer
- |
  stark
- |
  starkly
- |
  starkness
- |
  starless
- |
  starlet
- |
  starlight
- |
  starlike
- |
  starling
- |
  starlit
- |
  Starr
- |
  starred
- |
  starry
- |
  stars
- |
  start
- |
  starter
- |
  startle
- |
  startled
- |
  startling
- |
  startlingly
- |
  startup
- |
  starvation
- |
  starve
- |
  starveling
- |
  stash
- |
  stasis
- |
  state
- |
  statecraft
- |
  statehood
- |
  statehouse
- |
  stateless
- |
  stateliness
- |
  stately
- |
  statement
- |
  stateroom
- |
  States
- |
  stateside
- |
  statesman
- |
  stateswoman
- |
  statewide
- |
  static
- |
  statically
- |
  staticky
- |
  statics
- |
  station
- |
  stationary
- |
  stationer
- |
  stationery
- |
  statism
- |
  statist
- |
  statistic
- |
  statistical
- |
  statistician
- |
  statistics
- |
  stative
- |
  stats
- |
  statuary
- |
  statue
- |
  statuesque
- |
  statuette
- |
  stature
- |
  status
- |
  statute
- |
  statutorily
- |
  statutory
- |
  staunch
- |
  staunchly
- |
  staunchness
- |
  stave
- |
  staves
- |
  Stavropol
- |
  stays
- |
  stead
- |
  steadfast
- |
  steadfastly
- |
  steadily
- |
  steadiness
- |
  steady
- |
  steak
- |
  steal
- |
  stealer
- |
  stealth
- |
  stealthily
- |
  stealthiness
- |
  stealthy
- |
  steam
- |
  steamboat
- |
  steamer
- |
  steamfitter
- |
  steamfitting
- |
  steamily
- |
  steaminess
- |
  steamroll
- |
  steamroller
- |
  steamship
- |
  steamy
- |
  steatite
- |
  steed
- |
  steel
- |
  Steele
- |
  steeliness
- |
  steelworks
- |
  steely
- |
  steelyard
- |
  steep
- |
  steeped
- |
  steepen
- |
  steeple
- |
  steeplechase
- |
  steeplejack
- |
  steeply
- |
  steepness
- |
  steer
- |
  steerable
- |
  steerage
- |
  steerer
- |
  steering
- |
  steersman
- |
  Stefan
- |
  stegosaur
- |
  stegosaurus
- |
  Steichen
- |
  Stein
- |
  stein
- |
  Steinbeck
- |
  Steinem
- |
  stela
- |
  stelae
- |
  stele
- |
  Stella
- |
  stellar
- |
  stemless
- |
  stemma
- |
  stemmata
- |
  stemmatics
- |
  stemmed
- |
  stemware
- |
  stemwinder
- |
  stench
- |
  stencil
- |
  Stendhal
- |
  steno
- |
  stenographer
- |
  stenographic
- |
  stenography
- |
  stenosed
- |
  stenosing
- |
  stenosis
- |
  stenotic
- |
  stent
- |
  stentor
- |
  stentorian
- |
  stepbrother
- |
  stepchild
- |
  stepchildren
- |
  stepdaughter
- |
  stepfather
- |
  Stephan
- |
  Stephanie
- |
  Stephen
- |
  stepladder
- |
  stepmother
- |
  stepparent
- |
  steppe
- |
  stepper
- |
  stepsister
- |
  stepson
- |
  stere
- |
  stereo
- |
  stereograph
- |
  stereography
- |
  stereophonic
- |
  stereopticon
- |
  stereoscope
- |
  stereoscopic
- |
  stereoscopy
- |
  stereotype
- |
  stereotyped
- |
  stereotypic
- |
  sterile
- |
  sterilely
- |
  sterilise
- |
  sterility
- |
  sterilize
- |
  sterilizer
- |
  Sterling
- |
  sterling
- |
  Stern
- |
  stern
- |
  sterna
- |
  Sterne
- |
  sternly
- |
  sternness
- |
  sternum
- |
  sternutation
- |
  steroid
- |
  steroidal
- |
  sterol
- |
  stertorous
- |
  stertorously
- |
  stethoscope
- |
  stetson
- |
  Steuben
- |
  Steve
- |
  stevedore
- |
  Steven
- |
  Stevens
- |
  Stevenson
- |
  steward
- |
  stewardess
- |
  stewardship
- |
  Stewart
- |
  sthenic
- |
  stick
- |
  sticker
- |
  stickily
- |
  stickiness
- |
  stickleback
- |
  stickler
- |
  stickpin
- |
  sticks
- |
  stickup
- |
  sticky
- |
  stiff
- |
  stiffen
- |
  stiffener
- |
  stiffening
- |
  stiffish
- |
  stiffly
- |
  stiffness
- |
  stifle
- |
  stifling
- |
  stiflingly
- |
  stigma
- |
  stigmata
- |
  stigmatic
- |
  stigmatize
- |
  stile
- |
  stiletto
- |
  still
- |
  stillbirth
- |
  stillborn
- |
  stillness
- |
  stilt
- |
  stilted
- |
  stiltedly
- |
  stiltedness
- |
  Stilton
- |
  stilts
- |
  stimulant
- |
  stimulate
- |
  stimulating
- |
  stimulation
- |
  stimulative
- |
  stimulator
- |
  stimuli
- |
  stimulus
- |
  sting
- |
  stinger
- |
  stingily
- |
  stinginess
- |
  stinging
- |
  stingray
- |
  stingy
- |
  stink
- |
  stinkbug
- |
  stinker
- |
  stinking
- |
  stinky
- |
  stint
- |
  stinter
- |
  stinting
- |
  stipend
- |
  stipple
- |
  stippler
- |
  stippling
- |
  stipulate
- |
  stipulation
- |
  stipulator
- |
  Stirling
- |
  stirrer
- |
  stirring
- |
  stirringly
- |
  stirrup
- |
  stitch
- |
  stitcher
- |
  stitchery
- |
  stitches
- |
  stitching
- |
  stoat
- |
  stochastic
- |
  stock
- |
  stockade
- |
  stockbroker
- |
  stockbroking
- |
  stockholder
- |
  Stockholm
- |
  stockily
- |
  stockiness
- |
  stockinet
- |
  stockinette
- |
  stocking
- |
  stockist
- |
  stockpile
- |
  Stockport
- |
  stockroom
- |
  stocks
- |
  stocktaking
- |
  Stockton
- |
  stocky
- |
  stockyard
- |
  stodgily
- |
  stodginess
- |
  stodgy
- |
  stogie
- |
  stogy
- |
  Stoic
- |
  stoic
- |
  stoical
- |
  stoically
- |
  Stoicism
- |
  stoicism
- |
  stoke
- |
  stoked
- |
  stoker
- |
  stole
- |
  stolen
- |
  stolid
- |
  stolidity
- |
  stolidly
- |
  stolidness
- |
  stolon
- |
  stoma
- |
  stomach
- |
  stomachache
- |
  stomacher
- |
  stomachic
- |
  stomata
- |
  stomp
- |
  Stone
- |
  stone
- |
  stoned
- |
  Stonehenge
- |
  stonemason
- |
  stonewall
- |
  stoneware
- |
  stonewashed
- |
  stonework
- |
  stoney
- |
  stonily
- |
  stoniness
- |
  stony
- |
  stood
- |
  stooge
- |
  stool
- |
  stoop
- |
  stooping
- |
  stopcock
- |
  stopgap
- |
  stoplight
- |
  stopover
- |
  stoppage
- |
  Stoppard
- |
  stopper
- |
  stopple
- |
  stopwatch
- |
  storage
- |
  store
- |
  storefront
- |
  storehouse
- |
  storekeeper
- |
  storeroom
- |
  stores
- |
  storey
- |
  storied
- |
  stork
- |
  storm
- |
  stormily
- |
  storminess
- |
  storming
- |
  stormy
- |
  Stornoway
- |
  story
- |
  storyboard
- |
  storybook
- |
  storyline
- |
  storyteller
- |
  storytelling
- |
  stotinka
- |
  stoup
- |
  stout
- |
  stouthearted
- |
  stoutly
- |
  stoutness
- |
  stove
- |
  stovepipe
- |
  stowage
- |
  stowaway
- |
  Stowe
- |
  Strabane
- |
  strabismal
- |
  strabismic
- |
  strabismus
- |
  straddle
- |
  straddler
- |
  Stradivari
- |
  Stradivarius
- |
  strafe
- |
  strafer
- |
  straggle
- |
  straggler
- |
  straggly
- |
  straight
- |
  straightaway
- |
  straightedge
- |
  straighten
- |
  straightener
- |
  straightly
- |
  straightness
- |
  straightway
- |
  strain
- |
  strained
- |
  strainer
- |
  strains
- |
  strait
- |
  straiten
- |
  straitened
- |
  straitjacket
- |
  straitlaced
- |
  straitly
- |
  straitness
- |
  straits
- |
  strand
- |
  stranded
- |
  strange
- |
  strangely
- |
  strangeness
- |
  stranger
- |
  strangle
- |
  stranglehold
- |
  strangler
- |
  strangulate
- |
  strap
- |
  strapless
- |
  strappado
- |
  strapped
- |
  strapping
- |
  Strasbourg
- |
  strata
- |
  stratagem
- |
  strategic
- |
  strategical
- |
  strategics
- |
  strategist
- |
  strategy
- |
  Strathclyde
- |
  strati
- |
  stratified
- |
  stratify
- |
  stratigraphy
- |
  stratocracy
- |
  stratosphere
- |
  stratum
- |
  stratus
- |
  Strauss
- |
  Stravinsky
- |
  straw
- |
  strawberry
- |
  strawflower
- |
  stray
- |
  streak
- |
  streaker
- |
  streaky
- |
  stream
- |
  streambed
- |
  streamer
- |
  streamlet
- |
  streamline
- |
  streamlined
- |
  street
- |
  streetcar
- |
  streetlight
- |
  streetwalker
- |
  streetwise
- |
  strength
- |
  strengthen
- |
  strengthener
- |
  strenuous
- |
  strenuously
- |
  strep
- |
  streptococci
- |
  streptomycin
- |
  stress
- |
  stressed
- |
  stressful
- |
  stressor
- |
  stretch
- |
  stretchable
- |
  stretched
- |
  stretcher
- |
  stretching
- |
  stretchy
- |
  strew
- |
  strewn
- |
  stria
- |
  striae
- |
  striate
- |
  striated
- |
  striation
- |
  stricken
- |
  strict
- |
  strictly
- |
  strictness
- |
  stricture
- |
  strictured
- |
  stridden
- |
  stride
- |
  stridence
- |
  stridency
- |
  strident
- |
  stridently
- |
  strider
- |
  strides
- |
  stridor
- |
  stridulant
- |
  stridulate
- |
  stridulation
- |
  stridulatory
- |
  strife
- |
  strike
- |
  strikeout
- |
  striker
- |
  striking
- |
  strikingly
- |
  Strindberg
- |
  string
- |
  stringed
- |
  stringency
- |
  stringent
- |
  stringently
- |
  stringer
- |
  stringiness
- |
  strings
- |
  stringy
- |
  strip
- |
  stripe
- |
  striped
- |
  stripling
- |
  stripper
- |
  striptease
- |
  stripteaser
- |
  strive
- |
  striven
- |
  striving
- |
  strobe
- |
  stroboscope
- |
  stroboscopic
- |
  strode
- |
  stroke
- |
  stroll
- |
  stroller
- |
  Stromboli
- |
  strong
- |
  strongbox
- |
  stronghold
- |
  strongish
- |
  strongly
- |
  strongman
- |
  strongroom
- |
  strontium
- |
  strop
- |
  strophe
- |
  strophic
- |
  strove
- |
  struck
- |
  structural
- |
  structurally
- |
  structure
- |
  structured
- |
  strudel
- |
  struggle
- |
  struggler
- |
  strum
- |
  strumpet
- |
  strung
- |
  strut
- |
  strutter
- |
  struttingly
- |
  strychnine
- |
  Stuart
- |
  stubbiness
- |
  stubble
- |
  stubbly
- |
  stubborn
- |
  stubbornly
- |
  stubbornness
- |
  stubby
- |
  stucco
- |
  stuccoed
- |
  stuck
- |
  studbook
- |
  studded
- |
  studding
- |
  student
- |
  studentship
- |
  studied
- |
  studiedly
- |
  studies
- |
  studio
- |
  studious
- |
  studiously
- |
  studiousness
- |
  study
- |
  stuff
- |
  stuffed
- |
  stuffily
- |
  stuffiness
- |
  stuffing
- |
  stuffy
- |
  stultifier
- |
  stultify
- |
  stultifying
- |
  stumble
- |
  stumbler
- |
  stump
- |
  stumper
- |
  stumpy
- |
  stung
- |
  stunk
- |
  stunned
- |
  stunning
- |
  stunningly
- |
  stunt
- |
  stunted
- |
  stupa
- |
  stupefaction
- |
  stupefied
- |
  stupefier
- |
  stupefy
- |
  stupefying
- |
  stupefyingly
- |
  stupendous
- |
  stupendously
- |
  stupid
- |
  stupidity
- |
  stupidly
- |
  stupidness
- |
  stupor
- |
  stuporous
- |
  sturdily
- |
  sturdiness
- |
  sturdy
- |
  sturgeon
- |
  stutter
- |
  stutterer
- |
  stuttering
- |
  stutteringly
- |
  Stuttgart
- |
  Stuyvesant
- |
  Stygian
- |
  style
- |
  styli
- |
  styling
- |
  stylised
- |
  stylish
- |
  stylishly
- |
  stylishness
- |
  stylist
- |
  stylistic
- |
  stylistics
- |
  stylize
- |
  stylized
- |
  stylus
- |
  stymie
- |
  stymy
- |
  stypsis
- |
  styptic
- |
  styrene
- |
  Styrofoam
- |
  styrofoam
- |
  suasion
- |
  suasive
- |
  suave
- |
  suavely
- |
  suaveness
- |
  suavity
- |
  subabdominal
- |
  subacute
- |
  subagency
- |
  subagent
- |
  subalpine
- |
  subaltern
- |
  subapical
- |
  subapically
- |
  subaqueous
- |
  subarctic
- |
  subarea
- |
  subarid
- |
  subassembly
- |
  subatomic
- |
  subaverage
- |
  subaxillary
- |
  subbasement
- |
  subbranch
- |
  subcategory
- |
  subcellular
- |
  subchapter
- |
  subclass
- |
  subclassify
- |
  subclinical
- |
  subcommander
- |
  subcommittee
- |
  subcompact
- |
  subconscious
- |
  subcontinent
- |
  subcontract
- |
  subcouncil
- |
  subcranial
- |
  subcultural
- |
  subculture
- |
  subcutaneous
- |
  subdeacon
- |
  subdean
- |
  subdeb
- |
  subdirector
- |
  subdirectory
- |
  subdistrict
- |
  subdivide
- |
  subdivider
- |
  subdivision
- |
  subduct
- |
  subduction
- |
  subdue
- |
  subdued
- |
  subduer
- |
  subdural
- |
  subentry
- |
  subfamily
- |
  subfield
- |
  subfloor
- |
  subflooring
- |
  subfreezing
- |
  subgenre
- |
  subgenus
- |
  subglacial
- |
  subgroup
- |
  subhead
- |
  subheading
- |
  subhuman
- |
  subindex
- |
  subindustry
- |
  subjacency
- |
  subjacent
- |
  subject
- |
  subjection
- |
  subjective
- |
  subjectively
- |
  subjectivity
- |
  subjectless
- |
  subjoin
- |
  subjugate
- |
  subjugation
- |
  subjugator
- |
  subjunctive
- |
  subkingdom
- |
  sublease
- |
  sublet
- |
  sublethal
- |
  sublethally
- |
  sublimate
- |
  sublimation
- |
  sublime
- |
  sublimely
- |
  sublimeness
- |
  subliminal
- |
  subliminally
- |
  sublimity
- |
  subliterate
- |
  sublunary
- |
  submarginal
- |
  submarine
- |
  submariner
- |
  submember
- |
  submerge
- |
  submergence
- |
  submergible
- |
  submerse
- |
  submersible
- |
  submersion
- |
  subminiature
- |
  subminimal
- |
  subminimum
- |
  submission
- |
  submissive
- |
  submissively
- |
  submit
- |
  submittal
- |
  submolecular
- |
  subnormal
- |
  subnormality
- |
  subnotebook
- |
  suboceanic
- |
  subofficer
- |
  suboptimal
- |
  suborbital
- |
  suborder
- |
  subordinate
- |
  suborn
- |
  subornation
- |
  suborner
- |
  subpar
- |
  subparagraph
- |
  subparallel
- |
  subpena
- |
  subphylum
- |
  subplot
- |
  subpoena
- |
  subprincipal
- |
  subproblem
- |
  subprogram
- |
  subregion
- |
  subrogate
- |
  subrogation
- |
  subroutine
- |
  subsample
- |
  subscribe
- |
  subscriber
- |
  subscript
- |
  subscription
- |
  subsection
- |
  subsegment
- |
  subsense
- |
  subsequent
- |
  subsequently
- |
  subseries
- |
  subservience
- |
  subserviency
- |
  subservient
- |
  subset
- |
  subside
- |
  subsidence
- |
  subsidiarily
- |
  subsidiarity
- |
  subsidiary
- |
  subsidise
- |
  subsidize
- |
  subsidized
- |
  subsidizing
- |
  subsidy
- |
  subsist
- |
  subsistence
- |
  subsistent
- |
  subsoil
- |
  subsonic
- |
  subspecialty
- |
  subspecies
- |
  substage
- |
  substance
- |
  substandard
- |
  substantial
- |
  substantiate
- |
  substantival
- |
  substantive
- |
  substation
- |
  substitute
- |
  substitution
- |
  substrata
- |
  substrate
- |
  substratum
- |
  substructure
- |
  subsumable
- |
  subsume
- |
  subsumption
- |
  subsurface
- |
  subsystem
- |
  subteen
- |
  subtemperate
- |
  subtenancy
- |
  subtenant
- |
  subtend
- |
  subterfuge
- |
  subterranean
- |
  subtext
- |
  subtextual
- |
  subthreshold
- |
  subtile
- |
  subtitle
- |
  subtitled
- |
  subtitles
- |
  subtle
- |
  subtleness
- |
  subtlety
- |
  subtly
- |
  subtopic
- |
  subtotal
- |
  subtract
- |
  subtraction
- |
  subtrahend
- |
  subtreasury
- |
  subtribe
- |
  subtropic
- |
  subtropical
- |
  subtropics
- |
  subtype
- |
  subunit
- |
  suburb
- |
  suburban
- |
  suburbanite
- |
  suburbia
- |
  suburbs
- |
  subvariety
- |
  subvent
- |
  subvention
- |
  subversion
- |
  subversive
- |
  subversively
- |
  subvert
- |
  subverter
- |
  subvisible
- |
  subvocal
- |
  subway
- |
  subzero
- |
  succeed
- |
  succeeder
- |
  succeeding
- |
  success
- |
  successful
- |
  successfully
- |
  succession
- |
  successional
- |
  successive
- |
  successively
- |
  successor
- |
  succinct
- |
  succinctly
- |
  succinctness
- |
  succor
- |
  succorless
- |
  succors
- |
  succotash
- |
  Succoth
- |
  succour
- |
  succubi
- |
  succubus
- |
  succulence
- |
  succulency
- |
  succulent
- |
  succulently
- |
  succumb
- |
  suchlike
- |
  Suchow
- |
  sucker
- |
  suckle
- |
  suckling
- |
  Sucre
- |
  sucre
- |
  sucrose
- |
  suction
- |
  suctional
- |
  Sudan
- |
  Sudanese
- |
  Sudbury
- |
  sudden
- |
  suddenly
- |
  suddenness
- |
  Sudeten
- |
  Sudetenland
- |
  sudorific
- |
  sudsy
- |
  suede
- |
  Suellen
- |
  Suetonius
- |
  suffer
- |
  sufferable
- |
  sufferably
- |
  sufferance
- |
  sufferer
- |
  suffering
- |
  suffice
- |
  sufficiency
- |
  sufficient
- |
  sufficiently
- |
  suffix
- |
  suffixation
- |
  suffixion
- |
  suffocate
- |
  suffocating
- |
  suffocation
- |
  Suffolk
- |
  suffragan
- |
  suffrage
- |
  suffrages
- |
  suffragette
- |
  suffragism
- |
  suffragist
- |
  suffuse
- |
  suffusion
- |
  suffusive
- |
  Sufic
- |
  Sufism
- |
  sugar
- |
  sugarcane
- |
  sugarcoat
- |
  sugared
- |
  sugariness
- |
  sugarless
- |
  sugarplum
- |
  sugary
- |
  suggest
- |
  suggestible
- |
  suggestion
- |
  suggestive
- |
  suggestively
- |
  Suharto
- |
  suicidal
- |
  suicidally
- |
  suicide
- |
  suitability
- |
  suitable
- |
  suitableness
- |
  suitably
- |
  suitcase
- |
  suite
- |
  suited
- |
  suiting
- |
  suitor
- |
  Sukarno
- |
  sukiyaki
- |
  Sukkot
- |
  Sukkoth
- |
  Sulawesi
- |
  Suleiman
- |
  sulfa
- |
  sulfate
- |
  sulfide
- |
  sulfite
- |
  sulfonamide
- |
  sulfur
- |
  sulfuric
- |
  sulfurous
- |
  sulkily
- |
  sulkiness
- |
  sulky
- |
  Sulla
- |
  sullen
- |
  sullenly
- |
  sullenness
- |
  Sullivan
- |
  sully
- |
  sulphate
- |
  sulphur
- |
  sulphurous
- |
  sultan
- |
  sultana
- |
  sultanate
- |
  sultrily
- |
  sultriness
- |
  sultry
- |
  sumac
- |
  sumach
- |
  Sumatra
- |
  Sumatran
- |
  Sumer
- |
  Sumerian
- |
  Sumgait
- |
  summarily
- |
  summariness
- |
  summarise
- |
  summarize
- |
  summary
- |
  summation
- |
  summational
- |
  summative
- |
  summer
- |
  summerhouse
- |
  summertime
- |
  summery
- |
  summit
- |
  summitry
- |
  summon
- |
  summoner
- |
  summons
- |
  Sumner
- |
  sumptuary
- |
  sumptuosity
- |
  sumptuous
- |
  sumptuously
- |
  sunbaked
- |
  sunbath
- |
  sunbathe
- |
  sunbather
- |
  sunbathing
- |
  sunbeam
- |
  Sunbelt
- |
  sunblock
- |
  sunbonnet
- |
  sunburn
- |
  sunburned
- |
  sunburnt
- |
  sunburst
- |
  Sunchon
- |
  Sunda
- |
  sundae
- |
  Sunday
- |
  sunder
- |
  sunderance
- |
  Sunderland
- |
  sundial
- |
  sundown
- |
  sundries
- |
  sundry
- |
  sunfish
- |
  sunflower
- |
  sunglasses
- |
  sunken
- |
  sunlamp
- |
  sunless
- |
  sunlight
- |
  sunlit
- |
  Sunna
- |
  Sunnah
- |
  Sunni
- |
  sunnily
- |
  sunniness
- |
  Sunnite
- |
  sunny
- |
  Sunnyvale
- |
  sunrise
- |
  sunroof
- |
  sunscreen
- |
  sunset
- |
  sunshade
- |
  sunshine
- |
  sunshiny
- |
  sunspot
- |
  sunstroke
- |
  sunsuit
- |
  suntan
- |
  suntanned
- |
  sunup
- |
  super
- |
  superable
- |
  superagency
- |
  superannuate
- |
  superb
- |
  superblock
- |
  superbly
- |
  superbomb
- |
  superbug
- |
  supercargo
- |
  supercharge
- |
  supercharger
- |
  supercilious
- |
  supercity
- |
  superclean
- |
  superconduct
- |
  supercool
- |
  superego
- |
  supereminent
- |
  superficial
- |
  superficies
- |
  superfine
- |
  superfluity
- |
  superfluous
- |
  supergalaxy
- |
  supergiant
- |
  superheat
- |
  superheavy
- |
  superhero
- |
  superhighway
- |
  superhuman
- |
  superhumanly
- |
  superimpose
- |
  superintend
- |
  Superior
- |
  superior
- |
  superiority
- |
  superiorly
- |
  superlative
- |
  superlatives
- |
  superliner
- |
  superlunary
- |
  Superman
- |
  superman
- |
  supermarket
- |
  supermodel
- |
  supermom
- |
  supernal
- |
  supernally
- |
  supernatural
- |
  supernormal
- |
  supernova
- |
  supernovae
- |
  superpatriot
- |
  superposable
- |
  superpose
- |
  superpower
- |
  superpremium
- |
  superrich
- |
  superscribe
- |
  superscript
- |
  supersecret
- |
  supersede
- |
  supersession
- |
  supersize
- |
  supersized
- |
  supersmart
- |
  supersonic
- |
  superspy
- |
  superstar
- |
  superstate
- |
  superstition
- |
  superstore
- |
  superstratum
- |
  superstrong
- |
  supersubtle
- |
  supersystem
- |
  supertanker
- |
  superthin
- |
  supervene
- |
  supervenient
- |
  supervening
- |
  supervention
- |
  supervise
- |
  supervision
- |
  supervisor
- |
  supervisory
- |
  superwoman
- |
  supine
- |
  supinely
- |
  supineness
- |
  supper
- |
  supplant
- |
  supplanter
- |
  supple
- |
  supplely
- |
  supplement
- |
  supplemental
- |
  suppleness
- |
  suppliance
- |
  suppliant
- |
  suppliantly
- |
  supplicant
- |
  supplicate
- |
  supplication
- |
  supplicatory
- |
  supplier
- |
  supplies
- |
  supply
- |
  support
- |
  supportable
- |
  supporter
- |
  supportive
- |
  supportively
- |
  supposal
- |
  suppose
- |
  supposed
- |
  supposedly
- |
  supposing
- |
  supposition
- |
  suppositious
- |
  suppository
- |
  suppress
- |
  suppressant
- |
  suppressible
- |
  suppression
- |
  suppressive
- |
  suppressor
- |
  suppurate
- |
  suppuration
- |
  suppurative
- |
  supra
- |
  supremacist
- |
  supremacy
- |
  supreme
- |
  supremely
- |
  supremeness
- |
  supremo
- |
  Surabaja
- |
  Surabaya
- |
  surah
- |
  sural
- |
  Surat
- |
  surcease
- |
  surcharge
- |
  surcingle
- |
  surefire
- |
  surefooted
- |
  surely
- |
  sureness
- |
  surety
- |
  suretyship
- |
  surface
- |
  surfboard
- |
  surfeit
- |
  surfer
- |
  surficial
- |
  surficially
- |
  surfing
- |
  surge
- |
  surgeon
- |
  surgery
- |
  surgical
- |
  surgically
- |
  Surinam
- |
  Suriname
- |
  Surinamese
- |
  surlily
- |
  surliness
- |
  surly
- |
  surmise
- |
  surmount
- |
  surmountable
- |
  surmounter
- |
  surname
- |
  surpass
- |
  surpassable
- |
  surpassing
- |
  surpassingly
- |
  surplice
- |
  surplus
- |
  surprise
- |
  surprised
- |
  surprising
- |
  surprisingly
- |
  surprize
- |
  surreal
- |
  surrealism
- |
  surrealist
- |
  surrealistic
- |
  surreality
- |
  surreally
- |
  surrender
- |
  Surrey
- |
  surrey
- |
  surrogacy
- |
  surrogate
- |
  surround
- |
  surrounding
- |
  surroundings
- |
  surtax
- |
  surtout
- |
  surveillance
- |
  survey
- |
  surveying
- |
  surveyor
- |
  survivable
- |
  survival
- |
  survivalist
- |
  survive
- |
  survivor
- |
  Susan
- |
  Susanna
- |
  Susannah
- |
  Susanne
- |
  susceptible
- |
  susceptibly
- |
  sushi
- |
  Susie
- |
  suspect
- |
  suspend
- |
  suspended
- |
  suspender
- |
  suspenders
- |
  suspense
- |
  suspenseful
- |
  suspension
- |
  suspensory
- |
  suspicion
- |
  suspicious
- |
  suspiciously
- |
  suspiration
- |
  suspire
- |
  sustain
- |
  sustainable
- |
  sustainably
- |
  sustained
- |
  sustainedly
- |
  sustainer
- |
  sustaining
- |
  sustainment
- |
  sustenance
- |
  susurrant
- |
  susurrate
- |
  susurration
- |
  susurrous
- |
  susurrus
- |
  Sutherland
- |
  sutler
- |
  sutra
- |
  suttee
- |
  Sutton
- |
  suture
- |
  Suwon
- |
  Suzan
- |
  Suzann
- |
  Suzanne
- |
  suzerain
- |
  suzerainty
- |
  Suzhou
- |
  svelte
- |
  Svengali
- |
  Sverdlovsk
- |
  Swabia
- |
  Swabian
- |
  swaddle
- |
  swagged
- |
  swagger
- |
  Swahili
- |
  swain
- |
  swale
- |
  swallow
- |
  swallowtail
- |
  swami
- |
  swamp
- |
  swampiness
- |
  swampland
- |
  swampy
- |
  swank
- |
  swankily
- |
  swankiness
- |
  swanky
- |
  swansdown
- |
  Swansea
- |
  sward
- |
  swarded
- |
  swarm
- |
  swart
- |
  swarthily
- |
  swarthiness
- |
  swarthy
- |
  swash
- |
  swashbuckler
- |
  swastika
- |
  swatch
- |
  swath
- |
  swathe
- |
  swatter
- |
  swayback
- |
  swaybacked
- |
  Swazi
- |
  Swaziland
- |
  swear
- |
  swearer
- |
  swearword
- |
  sweat
- |
  sweatband
- |
  sweater
- |
  sweatiness
- |
  sweating
- |
  sweatpants
- |
  sweats
- |
  sweatshirt
- |
  sweatshop
- |
  sweaty
- |
  Swede
- |
  swede
- |
  Sweden
- |
  Swedenborg
- |
  Swedish
- |
  sweep
- |
  sweeper
- |
  sweeping
- |
  sweepingly
- |
  sweepings
- |
  sweepstake
- |
  sweepstakes
- |
  sweet
- |
  sweetbread
- |
  sweetbriar
- |
  sweetbrier
- |
  sweetcorn
- |
  sweeten
- |
  sweetener
- |
  sweetening
- |
  sweetheart
- |
  sweetie
- |
  sweetish
- |
  sweetly
- |
  sweetmeat
- |
  sweetness
- |
  sweets
- |
  swell
- |
  swellhead
- |
  swellheaded
- |
  swelling
- |
  swelter
- |
  sweltering
- |
  swelteringly
- |
  swept
- |
  sweptback
- |
  swerve
- |
  Swift
- |
  swift
- |
  swiftly
- |
  swiftness
- |
  swill
- |
  swimmer
- |
  swimming
- |
  swimmingly
- |
  swimsuit
- |
  Swinburne
- |
  swindle
- |
  swindler
- |
  Swindon
- |
  swine
- |
  swing
- |
  swinge
- |
  swinger
- |
  swinging
- |
  swinish
- |
  swipe
- |
  swirl
- |
  swirly
- |
  swish
- |
  Swiss
- |
  switch
- |
  switchback
- |
  switchblade
- |
  switchboard
- |
  switcher
- |
  switchman
- |
  Switzerland
- |
  swivel
- |
  swivet
- |
  swollen
- |
  swoon
- |
  swoop
- |
  sword
- |
  swordfish
- |
  swordplay
- |
  swordsman
- |
  swordtail
- |
  swore
- |
  sworn
- |
  swung
- |
  sybarite
- |
  sybaritic
- |
  sybaritism
- |
  Sybil
- |
  sycamore
- |
  sycophancy
- |
  sycophant
- |
  sycophantic
- |
  Sydney
- |
  syllabary
- |
  syllabi
- |
  syllabic
- |
  syllabically
- |
  syllabicate
- |
  syllabicity
- |
  syllabify
- |
  syllable
- |
  syllabus
- |
  syllepses
- |
  syllepsis
- |
  sylleptic
- |
  syllogism
- |
  syllogistic
- |
  sylph
- |
  sylphic
- |
  sylphlike
- |
  sylvan
- |
  Sylvester
- |
  Sylvia
- |
  symbioses
- |
  symbiosis
- |
  symbiotic
- |
  symbol
- |
  symbolic
- |
  symbolical
- |
  symbolically
- |
  symbolise
- |
  Symbolism
- |
  symbolism
- |
  symbolist
- |
  symbolize
- |
  symbology
- |
  symmetric
- |
  symmetrical
- |
  symmetrize
- |
  symmetry
- |
  sympathetic
- |
  sympathies
- |
  sympathise
- |
  sympathiser
- |
  sympathize
- |
  sympathizer
- |
  sympathy
- |
  symphonic
- |
  symphony
- |
  symposia
- |
  symposium
- |
  symptom
- |
  symptomatic
- |
  synagog
- |
  synagogal
- |
  synagogue
- |
  synapse
- |
  synaptic
- |
  synch
- |
  synchronic
- |
  synchronise
- |
  synchronism
- |
  synchronize
- |
  synchronizer
- |
  synchronous
- |
  synchrony
- |
  syncopal
- |
  syncopate
- |
  syncopation
- |
  syncopator
- |
  syncope
- |
  syncretic
- |
  syncretism
- |
  syncretist
- |
  syncretistic
- |
  syndicate
- |
  syndicated
- |
  syndication
- |
  syndicator
- |
  syndrome
- |
  syndromic
- |
  synecdoche
- |
  synecdochic
- |
  synergetic
- |
  synergic
- |
  synergism
- |
  synergist
- |
  synergistic
- |
  synergy
- |
  synfuel
- |
  Synge
- |
  synod
- |
  synodal
- |
  synodic
- |
  synodical
- |
  synodically
- |
  synonym
- |
  synonymic
- |
  synonymity
- |
  synonymous
- |
  synonymously
- |
  synonymy
- |
  synopses
- |
  synopsis
- |
  synopsize
- |
  synoptic
- |
  synoptical
- |
  synoptically
- |
  Synoptics
- |
  synovia
- |
  synovial
- |
  syntactic
- |
  syntactical
- |
  syntax
- |
  syntheses
- |
  synthesis
- |
  synthesise
- |
  synthesiser
- |
  synthesize
- |
  synthesizer
- |
  synthetic
- |
  synthetical
- |
  synthetics
- |
  syphilis
- |
  syphilitic
- |
  syphon
- |
  Syracuse
- |
  Syria
- |
  Syrian
- |
  syringe
- |
  syrup
- |
  syrupy
- |
  system
- |
  systematic
- |
  systematical
- |
  systematize
- |
  systemic
- |
  systemically
- |
  systemize
- |
  systole
- |
  systolic
- |
  syzygial
- |
  syzygy
- |
  Szczecin
- |
  Szechuan
- |
  Szechwan
- |
  Szeged
- |
  Tabasco
- |
  tabbouleh
- |
  tabby
- |
  Tabernacle
- |
  tabernacle
- |
  tabernacled
- |
  tabescent
- |
  Tabitha
- |
  tabla
- |
  tablature
- |
  table
- |
  tableau
- |
  tableaux
- |
  tablecloth
- |
  tableland
- |
  tablespoon
- |
  tablet
- |
  tabletop
- |
  tableware
- |
  tabloid
- |
  taboo
- |
  tabor
- |
  tabouleh
- |
  tabouli
- |
  tabour
- |
  Tabriz
- |
  tabular
- |
  tabularly
- |
  tabulate
- |
  tabulated
- |
  tabulation
- |
  tabulator
- |
  tabuli
- |
  tacet
- |
  tachometer
- |
  tachometry
- |
  tachycardia
- |
  tacit
- |
  tacitly
- |
  tacitness
- |
  taciturn
- |
  taciturnity
- |
  taciturnly
- |
  Tacitus
- |
  tacker
- |
  tackily
- |
  tackiness
- |
  tackle
- |
  tackler
- |
  tacky
- |
  Tacoma
- |
  taconite
- |
  tactful
- |
  tactfully
- |
  tactic
- |
  tactical
- |
  tactically
- |
  tactician
- |
  tactics
- |
  tactile
- |
  tactilely
- |
  tactility
- |
  tactless
- |
  tactlessly
- |
  tactlessness
- |
  tadpole
- |
  Tadzhik
- |
  Tadzhikistan
- |
  Taegu
- |
  Taejon
- |
  taffeta
- |
  taffrail
- |
  taffy
- |
  Tagalog
- |
  tagger
- |
  Tagore
- |
  Tagus
- |
  tahini
- |
  Tahiti
- |
  Tahitian
- |
  Tahoe
- |
  Taichung
- |
  taiga
- |
  Taihoku
- |
  tailback
- |
  tailcoat
- |
  tailed
- |
  tailgate
- |
  tailgater
- |
  tailgating
- |
  tailings
- |
  tailless
- |
  taillight
- |
  tailor
- |
  tailored
- |
  tailoring
- |
  tailpipe
- |
  tails
- |
  tailspin
- |
  tailwind
- |
  Tainan
- |
  Taine
- |
  Taino
- |
  taint
- |
  tainted
- |
  taintless
- |
  Taipei
- |
  Taiwan
- |
  Taiwanese
- |
  Taiyuan
- |
  Tajik
- |
  Tajikistan
- |
  Takakkaw
- |
  taken
- |
  takeoff
- |
  takeout
- |
  takeover
- |
  taker
- |
  taking
- |
  takings
- |
  Taklimakan
- |
  Talcahuano
- |
  talcum
- |
  talebearer
- |
  talebearing
- |
  talent
- |
  talented
- |
  taler
- |
  talesman
- |
  Taliban
- |
  talisman
- |
  talismanic
- |
  talkative
- |
  talkatively
- |
  talker
- |
  talkie
- |
  talks
- |
  talky
- |
  Tallahassee
- |
  tallboy
- |
  tallier
- |
  Tallin
- |
  Tallinn
- |
  tallish
- |
  tallness
- |
  tallow
- |
  tallowy
- |
  tally
- |
  tallyho
- |
  Talmud
- |
  Talmudic
- |
  Talmudical
- |
  Talmudist
- |
  talon
- |
  taloned
- |
  talus
- |
  tamable
- |
  tamale
- |
  Tamara
- |
  tamarack
- |
  tamari
- |
  tamarind
- |
  tamarisk
- |
  Tamaulipas
- |
  tambala
- |
  tambour
- |
  tambourine
- |
  tameable
- |
  tameless
- |
  tamely
- |
  tameness
- |
  tamer
- |
  Tamerlane
- |
  Tamil
- |
  Tammuz
- |
  Tammy
- |
  Tampa
- |
  Tampan
- |
  tamper
- |
  Tampere
- |
  tamperer
- |
  tampering
- |
  Tampico
- |
  tampon
- |
  tanager
- |
  Tananarive
- |
  tanbark
- |
  Tancred
- |
  tandem
- |
  tandoori
- |
  Taney
- |
  Tanganyika
- |
  Tanganyikan
- |
  tangelo
- |
  tangency
- |
  tangent
- |
  tangential
- |
  tangentially
- |
  tangerine
- |
  tangibility
- |
  tangible
- |
  tangibleness
- |
  tangibles
- |
  tangibly
- |
  Tangier
- |
  Tangiers
- |
  tanginess
- |
  tangle
- |
  tangled
- |
  tango
- |
  Tangshan
- |
  tangy
- |
  tankard
- |
  tanker
- |
  tankful
- |
  tanned
- |
  tanner
- |
  tannery
- |
  tannin
- |
  Tanoan
- |
  tansy
- |
  tantalise
- |
  tantalize
- |
  tantalizer
- |
  tantalizing
- |
  tantalum
- |
  Tantalus
- |
  tantamount
- |
  tantra
- |
  tantric
- |
  tantrum
- |
  Tanya
- |
  Tanzania
- |
  Tanzanian
- |
  Taoism
- |
  Taoist
- |
  Taoistic
- |
  taper
- |
  tapered
- |
  taperingly
- |
  tapestry
- |
  tapeworm
- |
  taping
- |
  tapioca
- |
  tapir
- |
  tapper
- |
  tappet
- |
  taproom
- |
  taproot
- |
  tapster
- |
  tarantella
- |
  Taranto
- |
  tarantula
- |
  tarantulae
- |
  Tarawa
- |
  tardily
- |
  tardiness
- |
  tardy
- |
  tares
- |
  target
- |
  tariff
- |
  Tarkington
- |
  Tarlac
- |
  tarmac
- |
  tarnish
- |
  tarnishable
- |
  tarnished
- |
  Tarot
- |
  tarot
- |
  tarpaper
- |
  tarpaulin
- |
  tarpon
- |
  tarragon
- |
  tarrier
- |
  tarry
- |
  Tarrytown
- |
  tarsal
- |
  tarsi
- |
  Tarsus
- |
  tarsus
- |
  tartan
- |
  Tartar
- |
  tartar
- |
  tartaric
- |
  Tartary
- |
  tartlet
- |
  tartly
- |
  tartness
- |
  Tarzan
- |
  Tashkent
- |
  taskbar
- |
  taskforce
- |
  taskmaster
- |
  taskmistress
- |
  Tasman
- |
  Tasmania
- |
  Tasmanian
- |
  tassel
- |
  tasseled
- |
  tastable
- |
  taste
- |
  tasteful
- |
  tastefully
- |
  tastefulness
- |
  tasteless
- |
  tastelessly
- |
  taster
- |
  tastily
- |
  tastiness
- |
  tasting
- |
  tasty
- |
  tatami
- |
  Tatar
- |
  tater
- |
  Tatiana
- |
  Tatra
- |
  Tatry
- |
  tatter
- |
  tattered
- |
  tatters
- |
  tattersail
- |
  tatting
- |
  tattle
- |
  tattler
- |
  tattletale
- |
  tattoo
- |
  tattooed
- |
  tattooer
- |
  tattooist
- |
  taught
- |
  taunt
- |
  taunter
- |
  tauntingly
- |
  Taunton
- |
  taupe
- |
  taurine
- |
  tauromachian
- |
  tauromachic
- |
  tauromachy
- |
  Taurus
- |
  tauten
- |
  tautly
- |
  tautness
- |
  tautologic
- |
  tautological
- |
  tautologist
- |
  tautologize
- |
  tautologous
- |
  tautology
- |
  tautomerism
- |
  tavern
- |
  taverna
- |
  tawdrily
- |
  tawdriness
- |
  tawdry
- |
  tawniness
- |
  tawny
- |
  taxable
- |
  taxation
- |
  taxer
- |
  taxicab
- |
  taxidermist
- |
  taxidermy
- |
  taximeter
- |
  taxing
- |
  taxon
- |
  taxonomic
- |
  taxonomical
- |
  taxonomist
- |
  taxonomize
- |
  taxonomy
- |
  taxpayer
- |
  taxpaying
- |
  taxying
- |
  Taylor
- |
  Tayside
- |
  Tbilisi
- |
  Tchaikovsky
- |
  teaberry
- |
  teach
- |
  teachability
- |
  teachable
- |
  teacher
- |
  teaching
- |
  teachings
- |
  teacup
- |
  teacupful
- |
  teakettle
- |
  teammate
- |
  teamster
- |
  teamwork
- |
  teapot
- |
  tearable
- |
  teardrop
- |
  tearer
- |
  tearful
- |
  tearfully
- |
  tearily
- |
  teariness
- |
  tearjerker
- |
  tearoom
- |
  tears
- |
  teary
- |
  tease
- |
  teasel
- |
  teaseler
- |
  teaser
- |
  teasing
- |
  teasingly
- |
  teaspoon
- |
  teaspoonful
- |
  teaspoonsful
- |
  Tebaldi
- |
  Tebet
- |
  technetium
- |
  technic
- |
  technical
- |
  technicality
- |
  technically
- |
  technician
- |
  Technicolor
- |
  technique
- |
  technocracy
- |
  technocrat
- |
  technocratic
- |
  technologist
- |
  technology
- |
  tectonic
- |
  tectonically
- |
  tectonics
- |
  Tecumseh
- |
  Teddy
- |
  teddy
- |
  tedious
- |
  tediously
- |
  tediousness
- |
  tedium
- |
  teeming
- |
  teemingly
- |
  teenage
- |
  teenaged
- |
  teenager
- |
  teens
- |
  teensy
- |
  teeny
- |
  teenybopper
- |
  teepee
- |
  teeter
- |
  teeth
- |
  teethe
- |
  teething
- |
  teetotal
- |
  teetotaler
- |
  teetotalism
- |
  teetotaller
- |
  Teflon
- |
  Tegucigalpa
- |
  Teheran
- |
  Tehran
- |
  tektite
- |
  telecast
- |
  telecaster
- |
  telecommute
- |
  telecommuter
- |
  telegenic
- |
  telegram
- |
  telegraph
- |
  telegrapher
- |
  telegraphic
- |
  telegraphist
- |
  telegraphy
- |
  telekinesis
- |
  telekinetic
- |
  telemarketer
- |
  telemeter
- |
  telemetric
- |
  telemetrical
- |
  telemetry
- |
  telepathic
- |
  telepathist
- |
  telepathy
- |
  telephone
- |
  telephoner
- |
  telephonic
- |
  telephony
- |
  telephoto
- |
  teleplay
- |
  teleprinter
- |
  TelePrompTer
- |
  teleprompter
- |
  telescope
- |
  telescopic
- |
  Telescopium
- |
  teletext
- |
  telethon
- |
  Teletype
- |
  televise
- |
  television
- |
  telex
- |
  telic
- |
  telicity
- |
  Teller
- |
  teller
- |
  telling
- |
  tellingly
- |
  telltale
- |
  tellurian
- |
  telluric
- |
  tellurium
- |
  telly
- |
  telnet
- |
  temblor
- |
  temerity
- |
  Tempe
- |
  tempeh
- |
  temper
- |
  tempera
- |
  temperament
- |
  temperance
- |
  temperate
- |
  temperately
- |
  temperature
- |
  tempered
- |
  tempest
- |
  tempestuous
- |
  tempi
- |
  template
- |
  temple
- |
  tempo
- |
  temporal
- |
  temporally
- |
  temporarily
- |
  temporary
- |
  temporize
- |
  temporizer
- |
  tempt
- |
  temptation
- |
  tempted
- |
  tempter
- |
  tempting
- |
  temptingly
- |
  temptress
- |
  tempura
- |
  tenability
- |
  tenable
- |
  tenableness
- |
  tenably
- |
  tenacious
- |
  tenaciously
- |
  tenacity
- |
  tenancy
- |
  tenant
- |
  tenantable
- |
  tenantless
- |
  tenantry
- |
  tendency
- |
  tendentious
- |
  tender
- |
  tenderer
- |
  tenderfeet
- |
  tenderfoot
- |
  tenderize
- |
  tenderizer
- |
  tenderloin
- |
  tenderly
- |
  tenderness
- |
  tendinitis
- |
  tendinous
- |
  tendon
- |
  tendonitis
- |
  tendril
- |
  tenebrous
- |
  tenement
- |
  tenet
- |
  tenfold
- |
  tenge
- |
  Tennessean
- |
  Tennessee
- |
  Tennesseean
- |
  tennis
- |
  Tennyson
- |
  Tennysonian
- |
  Tenochtitlan
- |
  tenon
- |
  tenoner
- |
  tenor
- |
  tenour
- |
  tenpenny
- |
  tenpin
- |
  tenpins
- |
  tense
- |
  tensely
- |
  tenseness
- |
  tensile
- |
  tensility
- |
  tension
- |
  tensity
- |
  tensive
- |
  tensor
- |
  tentacle
- |
  tentacled
- |
  tentacular
- |
  tentative
- |
  tentatively
- |
  tenterhook
- |
  tenth
- |
  tenthly
- |
  tenuity
- |
  tenuous
- |
  tenuously
- |
  tenuousness
- |
  tenure
- |
  tenured
- |
  teosinte
- |
  Teotihuacan
- |
  tepee
- |
  Tepic
- |
  tepid
- |
  tepidity
- |
  tepidly
- |
  tepidness
- |
  tequila
- |
  terabyte
- |
  teraflops
- |
  teratogen
- |
  teratogenic
- |
  teratologist
- |
  teratology
- |
  terbium
- |
  tercentenary
- |
  tercet
- |
  teredines
- |
  teredo
- |
  Terence
- |
  Teresa
- |
  Tereshkova
- |
  tergiversate
- |
  teriyaki
- |
  termagant
- |
  terminable
- |
  terminal
- |
  terminally
- |
  terminate
- |
  termination
- |
  terminative
- |
  terminator
- |
  termini
- |
  terminology
- |
  terminus
- |
  termite
- |
  termly
- |
  terms
- |
  ternary
- |
  Terpsichore
- |
  terrace
- |
  terraced
- |
  terracotta
- |
  terrain
- |
  Terrance
- |
  terrapin
- |
  terraria
- |
  terrarium
- |
  terrazzo
- |
  Terrell
- |
  Terrence
- |
  terrene
- |
  terrestrial
- |
  Terri
- |
  terrible
- |
  terribleness
- |
  terribly
- |
  terrier
- |
  terrific
- |
  terrifically
- |
  terrified
- |
  terrify
- |
  terrifying
- |
  terrifyingly
- |
  Terrill
- |
  territorial
- |
  Territory
- |
  territory
- |
  terror
- |
  terrorise
- |
  terrorism
- |
  terrorist
- |
  terroristic
- |
  terrorize
- |
  terrorizer
- |
  Terry
- |
  terry
- |
  terrycloth
- |
  terse
- |
  tersely
- |
  terseness
- |
  Tertiary
- |
  tertiary
- |
  Tesla
- |
  tesla
- |
  tesselate
- |
  tesselation
- |
  tessellate
- |
  tessellated
- |
  tessellation
- |
  tessera
- |
  tesserae
- |
  tesseral
- |
  tessitura
- |
  testable
- |
  Testament
- |
  testament
- |
  testamentary
- |
  testate
- |
  testator
- |
  testatrices
- |
  testatrix
- |
  tester
- |
  testes
- |
  testicle
- |
  testicular
- |
  testifier
- |
  testify
- |
  testily
- |
  testimonial
- |
  testimony
- |
  testiness
- |
  testing
- |
  testis
- |
  testosterone
- |
  testy
- |
  tetanal
- |
  tetanus
- |
  tetchy
- |
  tether
- |
  Teton
- |
  tetra
- |
  tetracycline
- |
  tetrahedra
- |
  tetrahedral
- |
  tetrahedron
- |
  tetralogy
- |
  tetrameter
- |
  Teuton
- |
  Teutonic
- |
  Tevet
- |
  Texan
- |
  Texas
- |
  textbook
- |
  textile
- |
  textiles
- |
  textual
- |
  textually
- |
  textural
- |
  texture
- |
  textured
- |
  Thackeray
- |
  Thaddeus
- |
  Thailand
- |
  Thailander
- |
  thalami
- |
  thalamic
- |
  thalamus
- |
  thalassic
- |
  Thales
- |
  Thalesian
- |
  thalidomide
- |
  thallium
- |
  thallophyte
- |
  Thames
- |
  Thana
- |
  thanatology
- |
  thane
- |
  thanedom
- |
  thank
- |
  thankful
- |
  thankfully
- |
  thankfulness
- |
  thankless
- |
  thanklessly
- |
  thanks
- |
  Thanksgiving
- |
  thanksgiving
- |
  Thant
- |
  thatch
- |
  thatched
- |
  Thatcher
- |
  thatcher
- |
  thatching
- |
  thaumaturge
- |
  thaumaturgic
- |
  thaumaturgy
- |
  theanthropic
- |
  thearchy
- |
  theater
- |
  theatre
- |
  theatrical
- |
  theatrically
- |
  theatricals
- |
  theatrics
- |
  Thebae
- |
  Theban
- |
  thebe
- |
  Thebes
- |
  theft
- |
  thegn
- |
  their
- |
  theirs
- |
  theism
- |
  theist
- |
  theistic
- |
  theistical
- |
  Thelma
- |
  thematic
- |
  thematically
- |
  theme
- |
  themselves
- |
  thence
- |
  thenceforth
- |
  Theocracy
- |
  theocracy
- |
  theocrat
- |
  theocratic
- |
  Theocritus
- |
  Theodora
- |
  Theodore
- |
  Theodoric
- |
  Theodosius
- |
  theologian
- |
  theological
- |
  theology
- |
  theorem
- |
  theorematic
- |
  theoretic
- |
  theoretical
- |
  theoretician
- |
  theorise
- |
  theorist
- |
  theorize
- |
  theorizer
- |
  theorizing
- |
  theory
- |
  theosopher
- |
  theosophic
- |
  theosophical
- |
  theosophist
- |
  theosophy
- |
  therapeutic
- |
  therapeutics
- |
  therapeutist
- |
  therapist
- |
  therapy
- |
  Theravada
- |
  there
- |
  thereabout
- |
  thereabouts
- |
  thereafter
- |
  thereat
- |
  thereby
- |
  therefor
- |
  therefore
- |
  therefrom
- |
  therein
- |
  thereinafter
- |
  thereof
- |
  thereon
- |
  Theresa
- |
  Therese
- |
  thereto
- |
  theretofore
- |
  thereunto
- |
  thereupon
- |
  therewith
- |
  therewithal
- |
  thermal
- |
  thermally
- |
  thermals
- |
  thermistor
- |
  thermocline
- |
  thermocouple
- |
  thermometer
- |
  thermometric
- |
  thermometry
- |
  Thermopylae
- |
  Thermos
- |
  thermos
- |
  thermosphere
- |
  thermostat
- |
  thermostatic
- |
  thesaural
- |
  thesauri
- |
  thesaurus
- |
  these
- |
  theses
- |
  Theseus
- |
  thesis
- |
  Thespian
- |
  thespian
- |
  Thespis
- |
  Thessalian
- |
  Thessalonian
- |
  Thessalonica
- |
  Thessalonike
- |
  Thessaloniki
- |
  Thessaly
- |
  theta
- |
  theurgic
- |
  theurgical
- |
  theurgist
- |
  theurgy
- |
  thewless
- |
  thews
- |
  thewy
- |
  thiamin
- |
  thiamine
- |
  thick
- |
  thicken
- |
  thickener
- |
  thickening
- |
  thicket
- |
  thickheaded
- |
  thickish
- |
  thickly
- |
  thickness
- |
  thickset
- |
  thief
- |
  thieve
- |
  thievery
- |
  thieves
- |
  thievish
- |
  thigh
- |
  thighbone
- |
  thimble
- |
  thimbleful
- |
  Thimbu
- |
  Thimphu
- |
  thine
- |
  thing
- |
  thingamajig
- |
  things
- |
  think
- |
  thinkable
- |
  thinker
- |
  thinking
- |
  thinly
- |
  thinner
- |
  thinness
- |
  thinnish
- |
  third
- |
  thirdly
- |
  thirst
- |
  thirstily
- |
  thirstiness
- |
  thirsty
- |
  thirteen
- |
  thirteenth
- |
  thirtieth
- |
  thirty
- |
  thistle
- |
  thistledown
- |
  thither
- |
  thitherward
- |
  thole
- |
  tholepin
- |
  Thomas
- |
  Thomism
- |
  Thompson
- |
  Thomson
- |
  thong
- |
  thoraces
- |
  thoracic
- |
  thorax
- |
  Thoreau
- |
  Thoreauvian
- |
  thorium
- |
  thorn
- |
  thornily
- |
  thorniness
- |
  thorny
- |
  thorough
- |
  Thoroughbred
- |
  thoroughbred
- |
  thoroughfare
- |
  thoroughly
- |
  thoroughness
- |
  thorp
- |
  Thorpe
- |
  those
- |
  though
- |
  thought
- |
  thoughtful
- |
  thoughtfully
- |
  thoughtless
- |
  Thousand
- |
  thousand
- |
  thousandfold
- |
  thousandth
- |
  Thrace
- |
  Thracia
- |
  Thracian
- |
  thraldom
- |
  thrall
- |
  thralldom
- |
  thrash
- |
  thrasher
- |
  thrashing
- |
  thread
- |
  threadbare
- |
  threader
- |
  thready
- |
  threat
- |
  threaten
- |
  threatened
- |
  threatening
- |
  three
- |
  threefold
- |
  threepence
- |
  threescore
- |
  threesome
- |
  threnodial
- |
  threnodic
- |
  threnodist
- |
  threnody
- |
  thresh
- |
  thresher
- |
  threshing
- |
  threshold
- |
  threw
- |
  thrice
- |
  thrift
- |
  thriftily
- |
  thriftiness
- |
  thriftless
- |
  thrifty
- |
  thrill
- |
  thrilled
- |
  thriller
- |
  thrilling
- |
  thrillingly
- |
  thrive
- |
  thriven
- |
  thriver
- |
  thriving
- |
  throat
- |
  throated
- |
  throatily
- |
  throatiness
- |
  throaty
- |
  throb
- |
  throbbingly
- |
  throe
- |
  throes
- |
  thrombi
- |
  thromboses
- |
  thrombosis
- |
  thrombotic
- |
  thrombus
- |
  throne
- |
  throng
- |
  thronged
- |
  throttle
- |
  throttler
- |
  through
- |
  throughout
- |
  throughput
- |
  throughway
- |
  throve
- |
  throw
- |
  throwaway
- |
  throwback
- |
  thrower
- |
  throwing
- |
  thrown
- |
  thrum
- |
  thrush
- |
  thrust
- |
  thruster
- |
  thrustor
- |
  thruway
- |
  Thuban
- |
  Thucydides
- |
  thudding
- |
  thuggery
- |
  thuggish
- |
  thulium
- |
  thumb
- |
  thumbnail
- |
  thumbprint
- |
  thumbscrew
- |
  thumbtack
- |
  thump
- |
  thumping
- |
  thunder
- |
  thunderbolt
- |
  thunderclap
- |
  thundercloud
- |
  thunderer
- |
  thunderhead
- |
  thunderous
- |
  thunderously
- |
  thunderstorm
- |
  Thurber
- |
  Thurman
- |
  Thurrock
- |
  Thursday
- |
  thwack
- |
  thwacker
- |
  thwart
- |
  thyme
- |
  thymine
- |
  thymosin
- |
  thymus
- |
  thyristor
- |
  thyroid
- |
  thyroidal
- |
  thyroxin
- |
  thyroxine
- |
  thyself
- |
  Tianjin
- |
  tiara
- |
  Tiber
- |
  Tiberian
- |
  Tiberis
- |
  Tiberius
- |
  Tibesti
- |
  Tibet
- |
  Tibetan
- |
  tibia
- |
  tibiae
- |
  tibial
- |
  tical
- |
  ticker
- |
  ticket
- |
  ticking
- |
  tickle
- |
  tickled
- |
  tickler
- |
  ticklish
- |
  ticklishly
- |
  ticklishness
- |
  tickly
- |
  ticktock
- |
  tidal
- |
  tidally
- |
  tidbit
- |
  tiddlywinks
- |
  tideland
- |
  tidelands
- |
  tidewater
- |
  tideway
- |
  tidily
- |
  tidiness
- |
  tidings
- |
  tieback
- |
  tiebreaker
- |
  Tientsin
- |
  tiepin
- |
  Tiepolo
- |
  tiered
- |
  Tiffany
- |
  Tiflis
- |
  tiger
- |
  tigerish
- |
  tight
- |
  tighten
- |
  tightener
- |
  tightening
- |
  tightfisted
- |
  tightfitting
- |
  tightlipped
- |
  tightly
- |
  tightness
- |
  tightrope
- |
  tights
- |
  tightwad
- |
  tigress
- |
  Tigris
- |
  Tijuana
- |
  Tilburg
- |
  tilde
- |
  tiler
- |
  tiling
- |
  tillable
- |
  tillage
- |
  tiller
- |
  Tillich
- |
  tilter
- |
  tilth
- |
  timbale
- |
  timber
- |
  timbered
- |
  timberland
- |
  timberline
- |
  timbre
- |
  timbrel
- |
  Timbuktu
- |
  timekeeper
- |
  timekeeping
- |
  timeless
- |
  timelessly
- |
  timelessness
- |
  timeline
- |
  timeliness
- |
  timely
- |
  timeout
- |
  timepiece
- |
  timer
- |
  times
- |
  timeserver
- |
  timeserving
- |
  timetable
- |
  timeworn
- |
  timid
- |
  timidity
- |
  timidly
- |
  timidness
- |
  timing
- |
  Timisoara
- |
  timocracy
- |
  timocratic
- |
  Timor
- |
  timorous
- |
  timorously
- |
  timorousness
- |
  Timothy
- |
  timothy
- |
  timpani
- |
  timpanist
- |
  tinct
- |
  tincture
- |
  tinder
- |
  tinderbox
- |
  tined
- |
  tinfoil
- |
  tinge
- |
  tinged
- |
  tingle
- |
  tingler
- |
  tingling
- |
  tingly
- |
  tininess
- |
  tinker
- |
  tinkerer
- |
  tinkering
- |
  tinkle
- |
  tinkly
- |
  tinned
- |
  tinnily
- |
  tinniness
- |
  tinnitus
- |
  tinny
- |
  tinplate
- |
  tinsel
- |
  tinseled
- |
  tinselled
- |
  tinsmith
- |
  tinter
- |
  Tintoretto
- |
  tintype
- |
  tinware
- |
  tipper
- |
  tippet
- |
  tipping
- |
  tipple
- |
  tippler
- |
  tipsily
- |
  tipsiness
- |
  tipster
- |
  tipsy
- |
  tiptoe
- |
  tiptop
- |
  tirade
- |
  tiramisu
- |
  Tirana
- |
  Tirane
- |
  tired
- |
  tiredly
- |
  tiredness
- |
  tireless
- |
  tirelessly
- |
  tirelessness
- |
  Tiresias
- |
  tiresome
- |
  tiresomely
- |
  tiresomeness
- |
  tiring
- |
  Tirol
- |
  Tirolean
- |
  Tirolese
- |
  Tishri
- |
  tissue
- |
  Titan
- |
  titan
- |
  Titanic
- |
  titanic
- |
  titanically
- |
  titanium
- |
  titbit
- |
  tithable
- |
  tithe
- |
  tither
- |
  Titian
- |
  titian
- |
  Titianesque
- |
  Titicaca
- |
  titillate
- |
  titillating
- |
  titillation
- |
  titivate
- |
  titivation
- |
  title
- |
  titled
- |
  titleholder
- |
  titlist
- |
  titmice
- |
  titmouse
- |
  Titograd
- |
  titrate
- |
  titration
- |
  titter
- |
  tittivate
- |
  tittle
- |
  titular
- |
  Titus
- |
  tizzy
- |
  Tlaxcala
- |
  Tlingit
- |
  tmeses
- |
  tmesis
- |
  toadstool
- |
  toady
- |
  toadyism
- |
  toast
- |
  toaster
- |
  toastmaster
- |
  toasty
- |
  tobacco
- |
  tobacconist
- |
  Tobago
- |
  Tobagonian
- |
  Tobias
- |
  Tobit
- |
  toboggan
- |
  tobogganer
- |
  tobogganing
- |
  tobogganist
- |
  toccata
- |
  Tocqueville
- |
  tocsin
- |
  today
- |
  toddle
- |
  toddler
- |
  toddy
- |
  toehold
- |
  toenail
- |
  toffee
- |
  toffy
- |
  togaed
- |
  together
- |
  togetherness
- |
  toggery
- |
  toggle
- |
  Togliatti
- |
  Togolese
- |
  toile
- |
  toiler
- |
  toilet
- |
  toiletries
- |
  toiletry
- |
  toilette
- |
  toilful
- |
  toils
- |
  toilsome
- |
  toilworn
- |
  Tokay
- |
  token
- |
  tokenism
- |
  Tokyo
- |
  Tokyoite
- |
  tolar
- |
  Toledo
- |
  tolerability
- |
  tolerable
- |
  tolerably
- |
  tolerance
- |
  tolerant
- |
  tolerantly
- |
  tolerate
- |
  toleration
- |
  Tolkien
- |
  tollbooth
- |
  tollgate
- |
  tollhouse
- |
  tollway
- |
  Tolstoi
- |
  Tolstoy
- |
  Tolstoyan
- |
  Toltec
- |
  Toltecan
- |
  Toluca
- |
  toluene
- |
  Tolyatti
- |
  tomahawk
- |
  tomato
- |
  tomboy
- |
  tomboyish
- |
  tombstone
- |
  tomcat
- |
  tomfoolery
- |
  Tommie
- |
  Tommy
- |
  tomogram
- |
  tomograph
- |
  tomographic
- |
  tomography
- |
  tomorrow
- |
  Tomsk
- |
  tomtit
- |
  tonal
- |
  tonality
- |
  tonally
- |
  tonearm
- |
  toneless
- |
  tonelessly
- |
  toner
- |
  Tonga
- |
  Tongan
- |
  tongs
- |
  tongue
- |
  tongued
- |
  tongueless
- |
  tongues
- |
  tonic
- |
  tonically
- |
  tonicity
- |
  tonight
- |
  Tonkin
- |
  Tonkinese
- |
  tonnage
- |
  tonne
- |
  tonsil
- |
  tonsillar
- |
  tonsillitic
- |
  tonsillitis
- |
  tonsorial
- |
  tonsure
- |
  tontine
- |
  Tonya
- |
  toolbar
- |
  toolmaker
- |
  toolmaking
- |
  tooter
- |
  tooth
- |
  toothache
- |
  toothbrush
- |
  toothed
- |
  toothily
- |
  toothless
- |
  toothpaste
- |
  toothpick
- |
  toothsome
- |
  toothsomely
- |
  toothy
- |
  tootle
- |
  topaz
- |
  topcoat
- |
  topdressing
- |
  Topeka
- |
  toper
- |
  topflight
- |
  topgallant
- |
  topiarian
- |
  topiarist
- |
  topiary
- |
  topic
- |
  topical
- |
  topicality
- |
  topically
- |
  topknot
- |
  topless
- |
  topmast
- |
  topmost
- |
  topnotch
- |
  topographer
- |
  topographic
- |
  topography
- |
  topological
- |
  topologist
- |
  topology
- |
  toponym
- |
  toponymic
- |
  topper
- |
  topping
- |
  topple
- |
  topsail
- |
  topside
- |
  topsides
- |
  topsoil
- |
  topspin
- |
  toque
- |
  Torah
- |
  torah
- |
  Torbay
- |
  torch
- |
  torchbearer
- |
  torchlight
- |
  toreador
- |
  torero
- |
  toreutic
- |
  toreutics
- |
  torii
- |
  Torino
- |
  torment
- |
  tormenter
- |
  tormentingly
- |
  tormentor
- |
  tornado
- |
  Toronto
- |
  Torontonian
- |
  torpedo
- |
  torpid
- |
  torpidity
- |
  torpidly
- |
  torpor
- |
  torporific
- |
  torque
- |
  Torquemada
- |
  torquey
- |
  Torrance
- |
  torrent
- |
  torrential
- |
  Torreon
- |
  Torres
- |
  torrid
- |
  torridity
- |
  torridly
- |
  torridness
- |
  torsi
- |
  torsion
- |
  torsional
- |
  torsionally
- |
  torsionless
- |
  torso
- |
  torte
- |
  tortellini
- |
  tortfeasor
- |
  tortilla
- |
  tortious
- |
  tortoise
- |
  Tortola
- |
  tortoni
- |
  Tortuga
- |
  tortuosity
- |
  tortuous
- |
  tortuously
- |
  tortuousness
- |
  torture
- |
  torturer
- |
  torturous
- |
  torturously
- |
  Toryism
- |
  Toscanini
- |
  tossup
- |
  total
- |
  totalisator
- |
  totalitarian
- |
  totality
- |
  totalizator
- |
  totalizer
- |
  totally
- |
  totem
- |
  totemic
- |
  totemism
- |
  totemist
- |
  totemistic
- |
  totter
- |
  tottery
- |
  toucan
- |
  touch
- |
  touchable
- |
  touchdown
- |
  touche
- |
  touched
- |
  touchily
- |
  touchiness
- |
  touching
- |
  touchingly
- |
  touchline
- |
  touchscreen
- |
  touchstone
- |
  touchy
- |
  tough
- |
  toughen
- |
  toughener
- |
  toughly
- |
  toughness
- |
  Toulon
- |
  Toulouse
- |
  toupee
- |
  tourism
- |
  tourist
- |
  touristy
- |
  tourmaline
- |
  tournament
- |
  tourney
- |
  tourniquet
- |
  Tours
- |
  tousle
- |
  tousled
- |
  touter
- |
  towage
- |
  toward
- |
  towards
- |
  towboat
- |
  towel
- |
  toweling
- |
  towelling
- |
  tower
- |
  towered
- |
  towering
- |
  toweringly
- |
  towhead
- |
  towheaded
- |
  towhee
- |
  towline
- |
  townhouse
- |
  townie
- |
  townsfolk
- |
  township
- |
  townsman
- |
  townspeople
- |
  townswoman
- |
  towny
- |
  towpath
- |
  towrope
- |
  toxemia
- |
  toxemic
- |
  toxic
- |
  toxically
- |
  toxicity
- |
  toxicologic
- |
  toxicologist
- |
  toxicology
- |
  toxics
- |
  toxin
- |
  Toyama
- |
  Toynbee
- |
  Toyonaka
- |
  trace
- |
  traceability
- |
  traceable
- |
  tracer
- |
  tracery
- |
  trachea
- |
  tracheae
- |
  tracheal
- |
  tracheotomy
- |
  tracing
- |
  track
- |
  trackable
- |
  trackage
- |
  trackball
- |
  tracker
- |
  tracking
- |
  trackless
- |
  tracksuit
- |
  tract
- |
  tractability
- |
  tractable
- |
  tractably
- |
  traction
- |
  tractional
- |
  tractive
- |
  tractor
- |
  Tracy
- |
  tradable
- |
  trade
- |
  tradeable
- |
  trademark
- |
  tradeoff
- |
  trader
- |
  tradesman
- |
  tradespeople
- |
  tradeswoman
- |
  trading
- |
  tradition
- |
  traditional
- |
  traditionary
- |
  traditionist
- |
  traduce
- |
  traducement
- |
  traducer
- |
  Trafalgar
- |
  traffic
- |
  trafficker
- |
  trafficking
- |
  tragedian
- |
  tragedienne
- |
  tragedy
- |
  tragic
- |
  tragical
- |
  tragically
- |
  tragicomedy
- |
  tragicomic
- |
  tragicomical
- |
  trail
- |
  trailblazer
- |
  trailblazing
- |
  trailer
- |
  train
- |
  trainable
- |
  trained
- |
  trainee
- |
  trainer
- |
  training
- |
  trainman
- |
  traipse
- |
  trait
- |
  traitor
- |
  traitorous
- |
  traitorously
- |
  Trajan
- |
  trajectory
- |
  trammel
- |
  trammeler
- |
  trammels
- |
  tramontane
- |
  tramp
- |
  tramper
- |
  trample
- |
  trampler
- |
  trampoline
- |
  trampoliner
- |
  trampolinist
- |
  trance
- |
  tranquil
- |
  tranquility
- |
  tranquilize
- |
  tranquilizer
- |
  tranquillity
- |
  tranquillize
- |
  tranquilly
- |
  transact
- |
  transaction
- |
  transactions
- |
  transactor
- |
  transaxle
- |
  transceiver
- |
  transcend
- |
  transcendent
- |
  transcribe
- |
  transcriber
- |
  transcript
- |
  transdermal
- |
  transducer
- |
  transept
- |
  transeptal
- |
  transfer
- |
  transferable
- |
  transferal
- |
  transference
- |
  transferrer
- |
  transfigure
- |
  transfix
- |
  transfixed
- |
  transfixion
- |
  transfixt
- |
  transform
- |
  transformer
- |
  transfuse
- |
  transfuser
- |
  transfusion
- |
  transgender
- |
  transgress
- |
  transgressor
- |
  tranship
- |
  transience
- |
  transiency
- |
  transient
- |
  transiently
- |
  transistor
- |
  transit
- |
  transition
- |
  transitional
- |
  transitive
- |
  transitively
- |
  transitivity
- |
  transitorily
- |
  transitory
- |
  translatable
- |
  translate
- |
  translation
- |
  translator
- |
  translucence
- |
  translucency
- |
  translucent
- |
  transmigrate
- |
  transmission
- |
  transmissive
- |
  transmit
- |
  transmittal
- |
  transmitter
- |
  transmogrify
- |
  transmontane
- |
  transmutable
- |
  transmutably
- |
  transmute
- |
  transmuter
- |
  transoceanic
- |
  transom
- |
  transomed
- |
  transonic
- |
  transpacific
- |
  transparency
- |
  transparent
- |
  transpire
- |
  transplant
- |
  transpolar
- |
  transponder
- |
  transport
- |
  transporter
- |
  transports
- |
  transposable
- |
  transposal
- |
  transpose
- |
  transposer
- |
  transsexual
- |
  transship
- |
  transuranic
- |
  transuranium
- |
  Transvaal
- |
  transversal
- |
  transverse
- |
  transversely
- |
  transvestism
- |
  transvestite
- |
  Transylvania
- |
  trapdoor
- |
  trapeze
- |
  trapezia
- |
  trapezium
- |
  trapezoid
- |
  trapezoidal
- |
  trapped
- |
  trapper
- |
  trappings
- |
  Trappist
- |
  traps
- |
  trapshooting
- |
  trash
- |
  trashy
- |
  trauma
- |
  traumata
- |
  traumatic
- |
  traumatise
- |
  traumatize
- |
  traumatized
- |
  travail
- |
  travails
- |
  travel
- |
  traveler
- |
  traveling
- |
  traveller
- |
  travelling
- |
  travelog
- |
  travelogue
- |
  travels
- |
  traversable
- |
  traversal
- |
  traverse
- |
  traverser
- |
  travertine
- |
  travesty
- |
  Travis
- |
  trawl
- |
  trawler
- |
  treacherous
- |
  treachery
- |
  treacle
- |
  treacly
- |
  tread
- |
  treader
- |
  treadle
- |
  treadmill
- |
  treason
- |
  treasonable
- |
  treasonous
- |
  treasurable
- |
  treasure
- |
  treasured
- |
  treasurer
- |
  Treasury
- |
  treasury
- |
  treat
- |
  treatable
- |
  treater
- |
  treatise
- |
  treatment
- |
  treaty
- |
  treble
- |
  trebling
- |
  trebly
- |
  trecento
- |
  treeless
- |
  treelike
- |
  treetop
- |
  trefoil
- |
  trekker
- |
  trekking
- |
  trellis
- |
  trellised
- |
  trematode
- |
  tremble
- |
  trembler
- |
  tremendous
- |
  tremendously
- |
  tremolo
- |
  tremor
- |
  tremulous
- |
  tremulously
- |
  trench
- |
  trenchancy
- |
  trenchant
- |
  trenchantly
- |
  trencher
- |
  trencherman
- |
  trend
- |
  trendily
- |
  trendiness
- |
  trendy
- |
  Trent
- |
  Trenton
- |
  Trentonian
- |
  trepan
- |
  trephination
- |
  trephine
- |
  trepidation
- |
  trespass
- |
  trespasser
- |
  tress
- |
  tressel
- |
  tresses
- |
  trestle
- |
  Trevithick
- |
  Trevor
- |
  Triad
- |
  triad
- |
  triadic
- |
  triage
- |
  trial
- |
  trials
- |
  triangle
- |
  triangular
- |
  triangularly
- |
  triangulate
- |
  Triangulum
- |
  Triassic
- |
  triathlete
- |
  triathlon
- |
  tribal
- |
  tribalism
- |
  tribally
- |
  tribe
- |
  tribesman
- |
  tribeswoman
- |
  tribulation
- |
  tribulations
- |
  tribunal
- |
  tribunary
- |
  tribunate
- |
  tribune
- |
  tribuneship
- |
  tributary
- |
  tribute
- |
  trice
- |
  triceps
- |
  triceratops
- |
  trichina
- |
  trichinae
- |
  trichinosis
- |
  trick
- |
  tricker
- |
  trickery
- |
  trickily
- |
  trickiness
- |
  trickle
- |
  trickster
- |
  tricky
- |
  tricolor
- |
  tricolored
- |
  tricorn
- |
  tricorne
- |
  tricot
- |
  tricycle
- |
  trident
- |
  tried
- |
  triennial
- |
  triennially
- |
  Trieste
- |
  trifle
- |
  trifler
- |
  trifling
- |
  triflingly
- |
  trifocal
- |
  trifocals
- |
  trifoliate
- |
  triforia
- |
  triforium
- |
  trigger
- |
  triggered
- |
  triglyceride
- |
  trigonometry
- |
  trike
- |
  trilateral
- |
  trilby
- |
  trill
- |
  trillion
- |
  trillionth
- |
  trillium
- |
  trilobite
- |
  trilogy
- |
  trimaran
- |
  trimester
- |
  trimestral
- |
  trimestrial
- |
  trimeter
- |
  trimetric
- |
  trimetrical
- |
  trimly
- |
  trimmer
- |
  trimming
- |
  trimmings
- |
  trimness
- |
  trimonthly
- |
  trine
- |
  Trinidad
- |
  Trinidadian
- |
  Trinitarian
- |
  Trinity
- |
  trinity
- |
  trinket
- |
  trinketry
- |
  tripartite
- |
  tripartitely
- |
  tripartition
- |
  tripe
- |
  triphammer
- |
  triple
- |
  triplet
- |
  triplex
- |
  triplicate
- |
  triplication
- |
  triply
- |
  tripod
- |
  tripodal
- |
  Tripoli
- |
  Tripolitan
- |
  tripper
- |
  triptych
- |
  trireme
- |
  trisect
- |
  trisection
- |
  trisector
- |
  Tristan
- |
  Tristram
- |
  trite
- |
  tritely
- |
  triteness
- |
  tritium
- |
  Triton
- |
  triton
- |
  triturate
- |
  triumph
- |
  triumphal
- |
  triumphant
- |
  triumphantly
- |
  triumvir
- |
  triumviral
- |
  triumvirate
- |
  triumviri
- |
  triune
- |
  triunity
- |
  trivalency
- |
  trivalent
- |
  Trivandrum
- |
  trivet
- |
  trivia
- |
  trivial
- |
  triviality
- |
  trivialize
- |
  trivially
- |
  trivium
- |
  triweekly
- |
  Trobriand
- |
  trochaic
- |
  troche
- |
  trochee
- |
  trodden
- |
  troglodyte
- |
  troglodytic
- |
  troglodytism
- |
  Troia
- |
  troika
- |
  Troja
- |
  Trojan
- |
  troll
- |
  troller
- |
  trolley
- |
  trolleybus
- |
  trollop
- |
  Trollope
- |
  trolly
- |
  trombone
- |
  trombonist
- |
  tromp
- |
  Trondheim
- |
  troop
- |
  trooper
- |
  troops
- |
  troopship
- |
  trope
- |
  trophic
- |
  trophy
- |
  tropic
- |
  tropical
- |
  tropically
- |
  tropics
- |
  tropism
- |
  troposphere
- |
  tropospheric
- |
  troth
- |
  Trotski
- |
  Trotsky
- |
  Trotskyism
- |
  Trotskyist
- |
  Trotskyite
- |
  trotter
- |
  troubadour
- |
  trouble
- |
  troubled
- |
  troublemaker
- |
  troubler
- |
  troubleshoot
- |
  troublesome
- |
  troublespot
- |
  troubling
- |
  troublous
- |
  trough
- |
  trounce
- |
  trouncer
- |
  troupe
- |
  trouper
- |
  trouser
- |
  trousers
- |
  trousseau
- |
  trousseaux
- |
  trout
- |
  trove
- |
  Trowbridge
- |
  trowel
- |
  truancy
- |
  truant
- |
  truce
- |
  truck
- |
  truckage
- |
  trucker
- |
  trucking
- |
  truckle
- |
  truckler
- |
  truckload
- |
  truculence
- |
  truculency
- |
  truculent
- |
  truculently
- |
  Trudeau
- |
  trudge
- |
  trudger
- |
  Trudy
- |
  truehearted
- |
  truelove
- |
  trueness
- |
  truffle
- |
  truism
- |
  truistic
- |
  Trujillo
- |
  truly
- |
  Truman
- |
  trump
- |
  trumpery
- |
  trumpet
- |
  trumpeter
- |
  trumps
- |
  truncate
- |
  truncated
- |
  truncation
- |
  truncheon
- |
  trundle
- |
  trundler
- |
  trunk
- |
  trunks
- |
  Truro
- |
  truss
- |
  trust
- |
  trusted
- |
  trustee
- |
  trusteeship
- |
  truster
- |
  trustful
- |
  trustfully
- |
  trustfulness
- |
  trustily
- |
  trustiness
- |
  trusting
- |
  trustingly
- |
  trustworthy
- |
  trusty
- |
  Truth
- |
  truth
- |
  truthful
- |
  truthfully
- |
  truthfulness
- |
  trying
- |
  tryingly
- |
  tryout
- |
  tryst
- |
  tryster
- |
  tsardom
- |
  tsarina
- |
  tsarism
- |
  tsarist
- |
  tsetse
- |
  Tshombe
- |
  Tsinan
- |
  Tsingtao
- |
  Tsitsihar
- |
  tsunami
- |
  Tsvetaeva
- |
  Tswana
- |
  tubal
- |
  tubbiness
- |
  tubby
- |
  tubed
- |
  tubeless
- |
  tuber
- |
  tubercle
- |
  tubercular
- |
  tuberculin
- |
  tuberculoses
- |
  tuberculosis
- |
  tuberculous
- |
  tuberose
- |
  tuberous
- |
  tubing
- |
  Tubman
- |
  tubular
- |
  tubule
- |
  Tucana
- |
  tucker
- |
  Tucson
- |
  Tucuman
- |
  Tudor
- |
  Tuesday
- |
  tufted
- |
  tufter
- |
  tufty
- |
  tugboat
- |
  tughrik
- |
  tugrik
- |
  tuition
- |
  tuitional
- |
  tuitionary
- |
  tularemia
- |
  tulip
- |
  tulle
- |
  Tulsa
- |
  Tulsan
- |
  tumble
- |
  tumbledown
- |
  tumbler
- |
  tumbleweed
- |
  tumbrel
- |
  tumbril
- |
  tumescence
- |
  tumescent
- |
  tumescently
- |
  tumid
- |
  tumidity
- |
  tumidly
- |
  tummy
- |
  tumor
- |
  tumorous
- |
  tumour
- |
  tumuli
- |
  tumult
- |
  tumultuous
- |
  tumultuously
- |
  tumulus
- |
  tunability
- |
  tunable
- |
  tundra
- |
  tuneable
- |
  tuneful
- |
  tunefully
- |
  tunefulness
- |
  tuneless
- |
  tunelessly
- |
  tunelessness
- |
  tuner
- |
  tuneup
- |
  tungsten
- |
  Tungusic
- |
  tunic
- |
  Tunis
- |
  Tunisia
- |
  Tunisian
- |
  tunnel
- |
  tunneler
- |
  tunneller
- |
  tunny
- |
  tupelo
- |
  Tupian
- |
  Tupperware
- |
  tuque
- |
  turban
- |
  turbaned
- |
  turbid
- |
  turbidity
- |
  turbidly
- |
  turbidness
- |
  turbine
- |
  turbo
- |
  turbocharge
- |
  turbocharger
- |
  turbofan
- |
  turbojet
- |
  turboprop
- |
  turbot
- |
  turbulence
- |
  turbulent
- |
  turbulently
- |
  tureen
- |
  turfy
- |
  Turgenev
- |
  turgescence
- |
  turgescent
- |
  turgid
- |
  turgidity
- |
  turgidly
- |
  turgidness
- |
  Turin
- |
  Turing
- |
  Turkestan
- |
  Turkey
- |
  turkey
- |
  Turkic
- |
  Turkish
- |
  Turkmen
- |
  Turkmenian
- |
  Turkmenistan
- |
  Turku
- |
  turmeric
- |
  turmoil
- |
  turnabout
- |
  turnaround
- |
  turnbuckle
- |
  turncoat
- |
  turndown
- |
  Turner
- |
  turner
- |
  turnery
- |
  turning
- |
  turnip
- |
  turnkey
- |
  turnoff
- |
  turnon
- |
  turnout
- |
  turnover
- |
  turnpike
- |
  turnstile
- |
  turntable
- |
  turpentine
- |
  turpitude
- |
  turquois
- |
  turquoise
- |
  turret
- |
  turreted
- |
  turtle
- |
  turtledove
- |
  turtleneck
- |
  turtlenecked
- |
  turves
- |
  Tuscaloosa
- |
  Tuscan
- |
  Tuscany
- |
  Tuscarora
- |
  tusked
- |
  tusker
- |
  tussle
- |
  tussock
- |
  tussocky
- |
  Tutankhamen
- |
  Tutankhaten
- |
  tutelage
- |
  tutelar
- |
  tutelary
- |
  tutor
- |
  tutorial
- |
  tutoring
- |
  tutorship
- |
  Tutsi
- |
  tutti
- |
  Tutuila
- |
  Tuvalu
- |
  Tuvaluan
- |
  tuxedo
- |
  Tuxtla
- |
  twaddle
- |
  twaddler
- |
  Twain
- |
  twain
- |
  twang
- |
  twangy
- |
  tweak
- |
  Tweed
- |
  tweed
- |
  tweedily
- |
  tweediness
- |
  tweeds
- |
  tweedy
- |
  tween
- |
  tweet
- |
  tweeter
- |
  tweeze
- |
  tweezers
- |
  twelfth
- |
  twelve
- |
  twelvefold
- |
  twelvemonth
- |
  twentieth
- |
  twenty
- |
  twerp
- |
  twice
- |
  twiddle
- |
  twiddler
- |
  twiddly
- |
  twiggy
- |
  twilight
- |
  twilit
- |
  twill
- |
  twilled
- |
  twine
- |
  twiner
- |
  twinge
- |
  twinight
- |
  twinkle
- |
  twinkler
- |
  twinkling
- |
  twinkly
- |
  twinning
- |
  twirl
- |
  twirler
- |
  twirly
- |
  twist
- |
  twisted
- |
  twister
- |
  twisty
- |
  twitch
- |
  twitchy
- |
  twitter
- |
  twittery
- |
  twixt
- |
  twofer
- |
  twofold
- |
  twohanded
- |
  twopence
- |
  twopenny
- |
  twosome
- |
  tychism
- |
  tycoon
- |
  tycoonery
- |
  tying
- |
  Tyler
- |
  tympana
- |
  tympani
- |
  tympanic
- |
  tympanist
- |
  tympanum
- |
  Tyndale
- |
  typecast
- |
  typeface
- |
  typescript
- |
  typeset
- |
  typesetter
- |
  typesetting
- |
  typewrite
- |
  typewriter
- |
  typewriting
- |
  typewritten
- |
  typewrote
- |
  typhoid
- |
  typhoon
- |
  typhous
- |
  typhus
- |
  typical
- |
  typicality
- |
  typically
- |
  typicalness
- |
  typification
- |
  typifier
- |
  typify
- |
  typing
- |
  typist
- |
  typographer
- |
  typographic
- |
  typography
- |
  typological
- |
  typologist
- |
  typology
- |
  tyrannic
- |
  tyrannical
- |
  tyrannically
- |
  tyrannicidal
- |
  tyrannicide
- |
  tyrannize
- |
  tyrannizer
- |
  tyrannosaur
- |
  tyrannous
- |
  tyrannously
- |
  tyranny
- |
  tyrant
- |
  Tyrian
- |
  Tyrol
- |
  Tyrolean
- |
  Tyrolese
- |
  Tyrone
- |
  Tyrrhenian
- |
  tzarina
- |
  Tzupo
- |
  Ubangi
- |
  Ubermensch
- |
  Ubermenschen
- |
  ubiety
- |
  ubiquitarian
- |
  ubiquitous
- |
  ubiquitously
- |
  ubiquity
- |
  Uccello
- |
  udder
- |
  Uffizi
- |
  ufologist
- |
  ufology
- |
  Uganda
- |
  Ugandan
- |
  uglification
- |
  uglify
- |
  ugliness
- |
  Ugric
- |
  ukase
- |
  ukelele
- |
  Ukraine
- |
  Ukrainian
- |
  ukulele
- |
  Ulaanbaatar
- |
  ulcer
- |
  ulcerate
- |
  ulceration
- |
  ulcerative
- |
  ulcerous
- |
  ullage
- |
  ulnae
- |
  ulnar
- |
  Ulsan
- |
  Ulster
- |
  ulster
- |
  ulterior
- |
  ultima
- |
  ultimacy
- |
  ultimata
- |
  ultimate
- |
  ultimately
- |
  ultimatum
- |
  ultimo
- |
  ultra
- |
  ultrafiche
- |
  ultrahigh
- |
  ultraliberal
- |
  ultralight
- |
  ultramarine
- |
  ultramodern
- |
  ultramontane
- |
  ultrapure
- |
  ultrashort
- |
  ultrasonic
- |
  ultrasonics
- |
  ultrasound
- |
  ultraviolet
- |
  ululate
- |
  ululation
- |
  Ulyanovsk
- |
  Ulysses
- |
  umbel
- |
  umbellate
- |
  umber
- |
  umbilical
- |
  umbilici
- |
  umbilicus
- |
  umbra
- |
  umbrae
- |
  umbrage
- |
  umbrageous
- |
  umbral
- |
  umbrella
- |
  Umbria
- |
  Umbrian
- |
  umbriferous
- |
  umiak
- |
  umlaut
- |
  umpire
- |
  umpteen
- |
  umpteenth
- |
  unabashed
- |
  unabated
- |
  unable
- |
  unabridged
- |
  unabsorbed
- |
  unabsorbent
- |
  unacademic
- |
  unaccented
- |
  unacceptable
- |
  unacceptably
- |
  unaccounted
- |
  unaccredited
- |
  unaccustomed
- |
  unachievable
- |
  unacquainted
- |
  unadapted
- |
  unaddressed
- |
  unadjusted
- |
  unadorned
- |
  unadvertised
- |
  unadvisable
- |
  unadvised
- |
  unadvisedly
- |
  unaesthetic
- |
  unaffected
- |
  unaffectedly
- |
  unaffiliated
- |
  unaffordable
- |
  unafraid
- |
  unaggressive
- |
  unaided
- |
  unalienable
- |
  unaligned
- |
  unalike
- |
  unallied
- |
  unallowable
- |
  unalloyed
- |
  unalloyedly
- |
  unalterable
- |
  unalterably
- |
  unaltered
- |
  unambiguous
- |
  unambitious
- |
  unanchored
- |
  unanimity
- |
  unanimous
- |
  unanimously
- |
  unannounced
- |
  unanswerable
- |
  unanswered
- |
  unapologetic
- |
  unapparent
- |
  unappealing
- |
  unappeasable
- |
  unappeased
- |
  unappetizing
- |
  unapproved
- |
  unarguable
- |
  unarguably
- |
  unarm
- |
  unarmed
- |
  unarmored
- |
  unartistic
- |
  unashamed
- |
  unashamedly
- |
  unasked
- |
  unassailable
- |
  unassertive
- |
  unassigned
- |
  unassisted
- |
  unassuming
- |
  unassumingly
- |
  unathletic
- |
  unattached
- |
  unattainable
- |
  unattempted
- |
  unattended
- |
  unattested
- |
  unattractive
- |
  unattributed
- |
  unauthentic
- |
  unauthorised
- |
  unauthorized
- |
  unavailable
- |
  unavailing
- |
  unavailingly
- |
  unavenged
- |
  unavoidable
- |
  unavoidably
- |
  unavowed
- |
  unawakened
- |
  unaware
- |
  unawareness
- |
  unawares
- |
  unbacked
- |
  unbaked
- |
  unbalanced
- |
  unbaptized
- |
  unbar
- |
  unbearable
- |
  unbearably
- |
  unbeatable
- |
  unbeaten
- |
  unbecoming
- |
  unbecomingly
- |
  unbefitting
- |
  unbeknown
- |
  unbeknownst
- |
  unbelief
- |
  unbelievable
- |
  unbelievably
- |
  unbeliever
- |
  unbelieving
- |
  unbeloved
- |
  unbend
- |
  unbending
- |
  unbendingly
- |
  unbent
- |
  unbiased
- |
  unbid
- |
  unbidden
- |
  unbind
- |
  unbleached
- |
  unblemished
- |
  unblenched
- |
  unblessed
- |
  unblest
- |
  unblinking
- |
  unblinkingly
- |
  unblock
- |
  unblushing
- |
  unblushingly
- |
  unbodied
- |
  unbolt
- |
  unbolted
- |
  unborn
- |
  unbosom
- |
  unbound
- |
  unbounded
- |
  unbowed
- |
  unbranched
- |
  unbranded
- |
  unbreakable
- |
  unbreathable
- |
  unbridgeable
- |
  unbridle
- |
  unbridled
- |
  unbroken
- |
  unbruised
- |
  unbrushed
- |
  unbuckle
- |
  unbudgeted
- |
  unbudging
- |
  unburden
- |
  unburied
- |
  unburned
- |
  unbutton
- |
  uncaged
- |
  uncanceled
- |
  uncannily
- |
  uncanniness
- |
  uncanny
- |
  uncanonical
- |
  uncap
- |
  uncaring
- |
  uncarpeted
- |
  uncashed
- |
  uncataloged
- |
  uncaught
- |
  unceasing
- |
  unceasingly
- |
  uncelebrated
- |
  uncensored
- |
  uncensured
- |
  uncertain
- |
  uncertainly
- |
  uncertainty
- |
  uncertified
- |
  unchain
- |
  unchallenged
- |
  unchangeable
- |
  unchangeably
- |
  unchanged
- |
  unchanging
- |
  unchaperoned
- |
  uncharged
- |
  uncharitable
- |
  uncharitably
- |
  uncharted
- |
  unchaste
- |
  unchastely
- |
  unchasteness
- |
  unchastity
- |
  unchecked
- |
  unchivalrous
- |
  unchristened
- |
  unchristian
- |
  unchurched
- |
  Uncial
- |
  uncial
- |
  uncirculated
- |
  uncivil
- |
  uncivilized
- |
  uncivilly
- |
  unclad
- |
  unclaimed
- |
  unclasp
- |
  unclassified
- |
  uncle
- |
  unclean
- |
  uncleaned
- |
  uncleanly
- |
  uncleanness
- |
  unclear
- |
  uncleared
- |
  unclench
- |
  uncloak
- |
  unclog
- |
  unclose
- |
  unclosed
- |
  unclothe
- |
  unclothed
- |
  unclouded
- |
  uncluttered
- |
  uncoated
- |
  uncoil
- |
  uncollected
- |
  uncolored
- |
  uncombed
- |
  uncombined
- |
  uncomely
- |
  uncomic
- |
  uncommercial
- |
  uncommitted
- |
  uncommon
- |
  uncommonly
- |
  uncommonness
- |
  uncompleted
- |
  uncompounded
- |
  unconcealed
- |
  unconcern
- |
  unconcerned
- |
  unconcluded
- |
  unconfined
- |
  unconfirmed
- |
  uncongenial
- |
  unconnected
- |
  unconquered
- |
  unconscious
- |
  unconsenting
- |
  unconsidered
- |
  unconsoled
- |
  unconsumed
- |
  uncontested
- |
  uncontrolled
- |
  unconverted
- |
  unconvinced
- |
  unconvincing
- |
  uncooked
- |
  uncork
- |
  uncorrected
- |
  uncorrupted
- |
  uncountable
- |
  uncounted
- |
  uncouple
- |
  uncourteous
- |
  uncouth
- |
  uncouthly
- |
  uncover
- |
  uncovered
- |
  uncrate
- |
  uncreative
- |
  uncredited
- |
  uncritical
- |
  uncritically
- |
  uncropped
- |
  uncross
- |
  uncrowded
- |
  uncrowned
- |
  unction
- |
  unctuous
- |
  unctuously
- |
  unctuousness
- |
  uncultivated
- |
  uncultured
- |
  uncured
- |
  uncurious
- |
  uncurl
- |
  uncurtained
- |
  uncustomary
- |
  uncut
- |
  undamaged
- |
  undamped
- |
  undated
- |
  undaunted
- |
  undauntedly
- |
  undebatable
- |
  undebatably
- |
  undeceivable
- |
  undeceivably
- |
  undeceive
- |
  undecided
- |
  undeclared
- |
  undecorated
- |
  undefeated
- |
  undefended
- |
  undefiled
- |
  undefinable
- |
  undefined
- |
  undemanding
- |
  undemocratic
- |
  undeniable
- |
  undeniably
- |
  undenied
- |
  undependable
- |
  under
- |
  underachieve
- |
  underact
- |
  underactive
- |
  underage
- |
  underaged
- |
  underarm
- |
  underbelly
- |
  underbid
- |
  underbidder
- |
  underbite
- |
  underbody
- |
  underbred
- |
  underbrush
- |
  undercharge
- |
  underclass
- |
  underclothes
- |
  undercoat
- |
  undercoating
- |
  undercover
- |
  undercroft
- |
  undercurrent
- |
  undercut
- |
  underdog
- |
  underdone
- |
  underdrawers
- |
  underdress
- |
  underexpose
- |
  underfed
- |
  underfeed
- |
  underfoot
- |
  underfur
- |
  undergarment
- |
  undergird
- |
  undergo
- |
  undergone
- |
  undergrad
- |
  underground
- |
  undergrowth
- |
  underhand
- |
  underhanded
- |
  underlain
- |
  underlay
- |
  underlie
- |
  underline
- |
  underling
- |
  underlip
- |
  underlying
- |
  undermine
- |
  underminer
- |
  undermost
- |
  underneath
- |
  underpaid
- |
  underpants
- |
  underpart
- |
  underpass
- |
  underpay
- |
  underpayment
- |
  underpin
- |
  underpinning
- |
  underplay
- |
  underproduce
- |
  underrate
- |
  underrated
- |
  underscore
- |
  undersea
- |
  underseas
- |
  undersell
- |
  undersexed
- |
  undershirt
- |
  undershoot
- |
  undershorts
- |
  undershot
- |
  underside
- |
  undersigned
- |
  undersize
- |
  undersized
- |
  underskirt
- |
  underslung
- |
  undersold
- |
  understaffed
- |
  understand
- |
  understate
- |
  understated
- |
  understood
- |
  understory
- |
  understudy
- |
  undersurface
- |
  undertake
- |
  undertaken
- |
  undertaker
- |
  undertaking
- |
  underthings
- |
  undertone
- |
  undertook
- |
  undertow
- |
  undertrick
- |
  undervalue
- |
  undervalued
- |
  underwater
- |
  underway
- |
  underwear
- |
  underweight
- |
  underwent
- |
  underwhelm
- |
  underworld
- |
  underwrite
- |
  underwriter
- |
  underwritten
- |
  underwrote
- |
  undeserved
- |
  undeservedly
- |
  undeserving
- |
  undesigned
- |
  undesigning
- |
  undesirable
- |
  undesirably
- |
  undesired
- |
  undetached
- |
  undetectable
- |
  undetected
- |
  undetermined
- |
  undeterred
- |
  undeveloped
- |
  undeviating
- |
  undiagnosed
- |
  undid
- |
  undies
- |
  undigested
- |
  undignified
- |
  undiluted
- |
  undiminished
- |
  undimmed
- |
  undine
- |
  undiplomatic
- |
  undirected
- |
  undiscerning
- |
  undisclosed
- |
  undiscovered
- |
  undisguised
- |
  undismayed
- |
  undisposed
- |
  undisputed
- |
  undissolved
- |
  undistressed
- |
  undisturbed
- |
  undivided
- |
  undocumented
- |
  undogmatic
- |
  undoing
- |
  undone
- |
  undoubled
- |
  undoubted
- |
  undoubtedly
- |
  undoubting
- |
  undramatic
- |
  undraped
- |
  undreamed
- |
  undreamt
- |
  undress
- |
  undressed
- |
  undrinkable
- |
  undue
- |
  undulant
- |
  undulate
- |
  undulately
- |
  undulating
- |
  undulation
- |
  undulatory
- |
  undulled
- |
  unduly
- |
  undutiful
- |
  undyed
- |
  undying
- |
  uneager
- |
  unearned
- |
  unearth
- |
  unearthly
- |
  unease
- |
  uneasily
- |
  uneasiness
- |
  uneasy
- |
  uneatable
- |
  uneaten
- |
  uneconomic
- |
  uneconomical
- |
  unedifying
- |
  unedited
- |
  uneducable
- |
  uneducated
- |
  unemotional
- |
  unemphatic
- |
  unemployable
- |
  unemployed
- |
  unemployment
- |
  unenclosed
- |
  unencumbered
- |
  unendangered
- |
  unending
- |
  unendorsed
- |
  unendurable
- |
  unendurably
- |
  unenforced
- |
  unenjoyable
- |
  unenriched
- |
  unenrolled
- |
  unentangled
- |
  unentered
- |
  unenviable
- |
  unequal
- |
  unequaled
- |
  unequalled
- |
  unequally
- |
  unequipped
- |
  unequivocal
- |
  unerring
- |
  unerringly
- |
  unescorted
- |
  unessential
- |
  unesthetic
- |
  unethical
- |
  unethically
- |
  uneven
- |
  unevenly
- |
  unevenness
- |
  uneventful
- |
  uneventfully
- |
  unexamined
- |
  unexampled
- |
  unexcelled
- |
  unexcited
- |
  unexciting
- |
  unexcused
- |
  unexercised
- |
  unexpected
- |
  unexpectedly
- |
  unexpended
- |
  unexpired
- |
  unexplained
- |
  unexplicit
- |
  unexploded
- |
  unexploited
- |
  unexplored
- |
  unexposed
- |
  unexpressed
- |
  unexpressive
- |
  unexpurgated
- |
  unfading
- |
  unfadingly
- |
  unfailing
- |
  unfailingly
- |
  unfair
- |
  unfairly
- |
  unfairness
- |
  unfaithful
- |
  unfaithfully
- |
  unfaltering
- |
  unfamiliar
- |
  unfamiliarly
- |
  unfasten
- |
  unfathomable
- |
  unfavorable
- |
  unfavorably
- |
  unfavourable
- |
  unfavourably
- |
  unfearing
- |
  unfeasible
- |
  unfed
- |
  unfederated
- |
  unfeeling
- |
  unfeelingly
- |
  unfeigned
- |
  unfelt
- |
  unfeminine
- |
  unfenced
- |
  unfermented
- |
  unfertilized
- |
  unfetter
- |
  unfettered
- |
  unfilial
- |
  unfilled
- |
  unfiltered
- |
  unfinished
- |
  unfit
- |
  unfitly
- |
  unfitness
- |
  unfitted
- |
  unfitting
- |
  unfittingly
- |
  unfix
- |
  unflagging
- |
  unflaggingly
- |
  unflappable
- |
  unflappably
- |
  unflattering
- |
  unflavored
- |
  unfledged
- |
  unflinching
- |
  unfocused
- |
  unfold
- |
  unfolded
- |
  unforced
- |
  unforeseen
- |
  unforetold
- |
  unforgivable
- |
  unforgiven
- |
  unforgiving
- |
  unforgotten
- |
  unformed
- |
  unformulated
- |
  unforsaken
- |
  unfortified
- |
  unfortunate
- |
  unfounded
- |
  unframed
- |
  unfree
- |
  unfreeze
- |
  unfrequented
- |
  unfriendly
- |
  unfrock
- |
  unfroze
- |
  unfrozen
- |
  unfruitful
- |
  unfulfilled
- |
  unfunded
- |
  unfunny
- |
  unfurl
- |
  unfurnished
- |
  unfussy
- |
  ungainliness
- |
  ungainly
- |
  Ungava
- |
  ungenerous
- |
  ungenerously
- |
  ungentle
- |
  ungerminated
- |
  unglamorous
- |
  unglazed
- |
  unglued
- |
  ungodliness
- |
  ungodly
- |
  ungovernable
- |
  ungoverned
- |
  ungraceful
- |
  ungracefully
- |
  ungracious
- |
  ungraciously
- |
  ungraded
- |
  ungrateful
- |
  ungratefully
- |
  ungratifying
- |
  unground
- |
  ungrounded
- |
  ungrudging
- |
  unguarded
- |
  unguent
- |
  unguided
- |
  ungulate
- |
  unhackneyed
- |
  unhallowed
- |
  unhampered
- |
  unhand
- |
  unhandsome
- |
  unhandy
- |
  unhappily
- |
  unhappiness
- |
  unhappy
- |
  unhardened
- |
  unharmed
- |
  unharmful
- |
  unharness
- |
  unharvested
- |
  unhatched
- |
  unhealed
- |
  unhealthful
- |
  unhealthily
- |
  unhealthy
- |
  unheard
- |
  unheated
- |
  unheeded
- |
  unheedful
- |
  unheedfully
- |
  unhelpful
- |
  unhelpfully
- |
  unheralded
- |
  unheroic
- |
  unhesitating
- |
  unhindered
- |
  unhinge
- |
  unhinged
- |
  unhistorical
- |
  unhitch
- |
  unholiness
- |
  unholy
- |
  unhonored
- |
  unhook
- |
  unhorse
- |
  unhoused
- |
  unhurried
- |
  unhurt
- |
  unhygienic
- |
  unhyphenated
- |
  unicameral
- |
  unicellular
- |
  unicorn
- |
  unicycle
- |
  unicyclist
- |
  unidentified
- |
  unidiomatic
- |
  unification
- |
  unified
- |
  uniform
- |
  uniformed
- |
  uniformity
- |
  uniformly
- |
  uniformness
- |
  unify
- |
  unilateral
- |
  unilaterally
- |
  unimaginable
- |
  unimaginably
- |
  unimpaired
- |
  unimpeded
- |
  unimportance
- |
  unimportant
- |
  unimposing
- |
  unimpressed
- |
  unimpressive
- |
  unimproved
- |
  uninfected
- |
  uninflected
- |
  uninfluenced
- |
  uninformed
- |
  uninhabited
- |
  uninhibited
- |
  uninitiated
- |
  uninjured
- |
  uninspired
- |
  uninspiring
- |
  uninstructed
- |
  uninsurable
- |
  uninsured
- |
  unintended
- |
  uninterested
- |
  uninvested
- |
  uninvited
- |
  uninviting
- |
  uninvitingly
- |
  uninvolved
- |
  Union
- |
  union
- |
  Unionism
- |
  unionism
- |
  unionist
- |
  unionization
- |
  unionize
- |
  unionized
- |
  unionizer
- |
  unique
- |
  uniquely
- |
  uniqueness
- |
  unironed
- |
  unisex
- |
  unisexual
- |
  unison
- |
  Unitarian
- |
  Unitarianism
- |
  unitarily
- |
  unitary
- |
  unite
- |
  united
- |
  unitize
- |
  unity
- |
  univalent
- |
  univalve
- |
  universal
- |
  Universalism
- |
  universalism
- |
  Universalist
- |
  universalist
- |
  universality
- |
  universalize
- |
  universally
- |
  universe
- |
  university
- |
  unjointed
- |
  unjust
- |
  unjustified
- |
  unjustly
- |
  unkempt
- |
  unkemptly
- |
  unkemptness
- |
  unkept
- |
  unkind
- |
  unkindliness
- |
  unkindly
- |
  unkindness
- |
  unkissed
- |
  unknowable
- |
  unknowing
- |
  unknowingly
- |
  unknown
- |
  unlabeled
- |
  unlace
- |
  unlade
- |
  unladen
- |
  unladylike
- |
  unlamented
- |
  unlatch
- |
  unlawful
- |
  unlawfully
- |
  unlawfulness
- |
  unleaded
- |
  unlearn
- |
  unlearned
- |
  unlearnedly
- |
  unleash
- |
  unleavened
- |
  unless
- |
  unlettered
- |
  unlicensed
- |
  unlighted
- |
  unlikable
- |
  unlike
- |
  unlikelihood
- |
  unlikeliness
- |
  unlikely
- |
  unlikeness
- |
  unlimber
- |
  unlimited
- |
  unlined
- |
  unlink
- |
  unlisted
- |
  unlit
- |
  unliterary
- |
  unlivable
- |
  unload
- |
  unloader
- |
  unlock
- |
  unloose
- |
  unloosen
- |
  unlovable
- |
  unloved
- |
  unlovely
- |
  unloving
- |
  unluckily
- |
  unluckiness
- |
  unlucky
- |
  unmade
- |
  unmagnified
- |
  unmake
- |
  unmalicious
- |
  unman
- |
  unmanageable
- |
  unmanageably
- |
  unmanly
- |
  unmanned
- |
  unmannered
- |
  unmanneredly
- |
  unmannerly
- |
  unmapped
- |
  unmarked
- |
  unmarketable
- |
  unmarred
- |
  unmarried
- |
  unmasculine
- |
  unmask
- |
  unmastered
- |
  unmatched
- |
  unmeaning
- |
  unmeant
- |
  unmeasurable
- |
  unmeasured
- |
  unmediated
- |
  unmeet
- |
  unmelodious
- |
  unmelted
- |
  unmemorized
- |
  unmended
- |
  unmentioned
- |
  unmerciful
- |
  unmercifully
- |
  unmerited
- |
  unmethodical
- |
  unmilitary
- |
  unmilled
- |
  unmindful
- |
  unmistakable
- |
  unmistakably
- |
  unmistaken
- |
  unmitigated
- |
  unmixed
- |
  unmodified
- |
  unmolded
- |
  unmolested
- |
  unmoor
- |
  unmoral
- |
  unmorality
- |
  unmotivated
- |
  unmounted
- |
  unmourned
- |
  unmovable
- |
  unmoved
- |
  unmown
- |
  unmuffle
- |
  unmusical
- |
  unmusically
- |
  unmuzzle
- |
  unmyelinated
- |
  unnameable
- |
  unnamed
- |
  unnatural
- |
  unnaturally
- |
  unnavigable
- |
  unnecessary
- |
  unneeded
- |
  unnegotiable
- |
  unneighborly
- |
  unnerve
- |
  unnerving
- |
  unnervingly
- |
  unnewsworthy
- |
  unnilhexium
- |
  unnilpentium
- |
  unnilquadium
- |
  unnoticeable
- |
  unnoticeably
- |
  unnoticed
- |
  unnumbered
- |
  unobliging
- |
  unobservant
- |
  unobserved
- |
  unobserving
- |
  unobstructed
- |
  unobtainable
- |
  unobtrusive
- |
  unoccupied
- |
  unoffended
- |
  unoffending
- |
  unoffensive
- |
  unoffered
- |
  unofficial
- |
  unofficially
- |
  unopened
- |
  unopposed
- |
  unordained
- |
  unorganized
- |
  unoriginal
- |
  unornament
- |
  unornamented
- |
  unorthodox
- |
  unorthodoxy
- |
  unowned
- |
  unpack
- |
  unpaged
- |
  unpaginated
- |
  unpaid
- |
  unpainted
- |
  unpaired
- |
  unpalatable
- |
  unpalatably
- |
  unparalleled
- |
  unpardonable
- |
  unpardonably
- |
  unpatented
- |
  unpatriotic
- |
  unpaved
- |
  unpeeled
- |
  unpeg
- |
  unpeople
- |
  unpeopled
- |
  unperceived
- |
  unperceptive
- |
  unperfected
- |
  unperformed
- |
  unperson
- |
  unpersuaded
- |
  unpersuasive
- |
  unperturbed
- |
  unpicked
- |
  unpile
- |
  unpin
- |
  unplanned
- |
  unplanted
- |
  unplayable
- |
  unplayed
- |
  unpleasant
- |
  unpleasantly
- |
  unpleased
- |
  unpleasing
- |
  unplowed
- |
  unplug
- |
  unplugged
- |
  unplumbed
- |
  unpoetic
- |
  unpoised
- |
  unpolished
- |
  unpolitical
- |
  unpolled
- |
  unpolluted
- |
  unpopular
- |
  unpopularity
- |
  unpopulated
- |
  unposed
- |
  unpractical
- |
  unpracticed
- |
  unpractised
- |
  unpredicted
- |
  unprejudiced
- |
  unprepared
- |
  unpreparedly
- |
  unpreserved
- |
  unpressed
- |
  unpretending
- |
  unpretty
- |
  unpriced
- |
  unprincipled
- |
  unprintable
- |
  unprivileged
- |
  unprocessed
- |
  unproclaimed
- |
  unproductive
- |
  unprofessed
- |
  unprofitable
- |
  unprofitably
- |
  unprogrammed
- |
  unprohibited
- |
  unpromising
- |
  unprompted
- |
  unpronounced
- |
  unpropitious
- |
  unprotected
- |
  unprotesting
- |
  unprovable
- |
  unproved
- |
  unproven
- |
  unprovided
- |
  unprovoked
- |
  unpublished
- |
  unpunished
- |
  unpurified
- |
  unqualified
- |
  unquenchable
- |
  unquenchably
- |
  unquenched
- |
  unquestioned
- |
  unquiet
- |
  unquotable
- |
  unquote
- |
  unraised
- |
  unrated
- |
  unratified
- |
  unravel
- |
  unreachable
- |
  unread
- |
  unreadable
- |
  unreadily
- |
  unreadiness
- |
  unready
- |
  unreal
- |
  unrealistic
- |
  unreality
- |
  unrealizable
- |
  unrealized
- |
  unreason
- |
  unreasonable
- |
  unreasonably
- |
  unreasoned
- |
  unreasoning
- |
  unreceptive
- |
  unreclaimed
- |
  unrecognized
- |
  unreconciled
- |
  unrecorded
- |
  unredeemable
- |
  unredeemed
- |
  unreel
- |
  unrefined
- |
  unreflecting
- |
  unreflective
- |
  unreformed
- |
  unregenerate
- |
  unregimented
- |
  unregistered
- |
  unregulated
- |
  unrehearsed
- |
  unrelated
- |
  unrelenting
- |
  unreliable
- |
  unreliably
- |
  unrelieved
- |
  unreligious
- |
  unremarkable
- |
  unremarkably
- |
  unremarked
- |
  unremembered
- |
  unremitting
- |
  unremorseful
- |
  unremovable
- |
  unremoved
- |
  unrenewed
- |
  unrented
- |
  unrepaid
- |
  unrepealed
- |
  unrepentant
- |
  unrepenting
- |
  unreported
- |
  unrepressed
- |
  unreproved
- |
  unrequited
- |
  unrequitedly
- |
  unresentful
- |
  unreserved
- |
  unreservedly
- |
  unresigned
- |
  unresistant
- |
  unresisting
- |
  unresolved
- |
  unrespectful
- |
  unresponsive
- |
  unrest
- |
  unrestful
- |
  unrestrained
- |
  unrestraint
- |
  unrestricted
- |
  unreturnable
- |
  unreturned
- |
  unrevealed
- |
  unrevenged
- |
  unrevised
- |
  unrevoked
- |
  unrewarded
- |
  unrewarding
- |
  unrhymed
- |
  unrhythmic
- |
  unriddle
- |
  unrighteous
- |
  unripe
- |
  unripened
- |
  unripeness
- |
  unrivaled
- |
  unrivalled
- |
  unrobe
- |
  unroll
- |
  unromantic
- |
  unroof
- |
  unruffled
- |
  unruliness
- |
  unruly
- |
  unsaddle
- |
  unsafe
- |
  unsafely
- |
  unsaid
- |
  unsalability
- |
  unsalable
- |
  unsalted
- |
  unsanctioned
- |
  unsanitary
- |
  unsatisfied
- |
  unsatisfying
- |
  unsaturate
- |
  unsaturated
- |
  unsaved
- |
  unsavorily
- |
  unsavoriness
- |
  unsavory
- |
  unsavoury
- |
  unsay
- |
  unscarred
- |
  unscathed
- |
  unscented
- |
  unscheduled
- |
  unscholarly
- |
  unschooled
- |
  unscientific
- |
  unscramble
- |
  unscratched
- |
  unscrew
- |
  unscripted
- |
  unscrupulous
- |
  unseal
- |
  unsealed
- |
  unsearchable
- |
  unseasonable
- |
  unseasonably
- |
  unseasoned
- |
  unseat
- |
  unseaworthy
- |
  unsecured
- |
  unseeded
- |
  unseeing
- |
  unseeingly
- |
  unseemliness
- |
  unseemly
- |
  unseen
- |
  unsegmented
- |
  unsegregated
- |
  unselfish
- |
  unselfishly
- |
  unsensitive
- |
  unsent
- |
  unserious
- |
  unsettle
- |
  unsettled
- |
  unsettling
- |
  unsettlingly
- |
  unsexual
- |
  unshackle
- |
  unshaded
- |
  unshakable
- |
  unshakably
- |
  unshaken
- |
  unshaped
- |
  unshapely
- |
  unshared
- |
  unshaved
- |
  unshaven
- |
  unsheathe
- |
  unshelled
- |
  unsheltered
- |
  unshielded
- |
  unship
- |
  unshockable
- |
  unshod
- |
  unshorn
- |
  unshrinking
- |
  unsifted
- |
  unsighted
- |
  unsightly
- |
  unsigned
- |
  unsinkable
- |
  unskilled
- |
  unskillful
- |
  unskillfully
- |
  unsliced
- |
  unsling
- |
  unslung
- |
  unsmiling
- |
  unsnap
- |
  unsnarl
- |
  unsociable
- |
  unsociably
- |
  unsocial
- |
  unsocially
- |
  unsoiled
- |
  unsold
- |
  unsoldierly
- |
  unsolicited
- |
  unsolvable
- |
  unsolved
- |
  unsorted
- |
  unsought
- |
  unsound
- |
  unsoundly
- |
  unsoundness
- |
  unsparing
- |
  unsparingly
- |
  unspeakable
- |
  unspeakably
- |
  unspecific
- |
  unspecified
- |
  unspent
- |
  unspiritual
- |
  unspoiled
- |
  unspoken
- |
  unspotted
- |
  unsprung
- |
  unstable
- |
  unstableness
- |
  unstably
- |
  unstained
- |
  unstamped
- |
  unstated
- |
  unsteadily
- |
  unsteadiness
- |
  unsteady
- |
  unsterile
- |
  unstick
- |
  unstinting
- |
  unstintingly
- |
  unstop
- |
  unstoppable
- |
  unstrap
- |
  unstressed
- |
  unstring
- |
  unstructured
- |
  unstrung
- |
  unstuck
- |
  unstudied
- |
  unstylish
- |
  unsubdued
- |
  unsubtle
- |
  unsuccess
- |
  unsuccessful
- |
  unsuitable
- |
  unsuitably
- |
  unsuited
- |
  unsullied
- |
  unsung
- |
  unsupervised
- |
  unsupported
- |
  unsuppressed
- |
  unsure
- |
  unsurely
- |
  unsureness
- |
  unsurpassed
- |
  unsurprised
- |
  unsurprising
- |
  unsuspected
- |
  unsuspecting
- |
  unsuspicious
- |
  unsustained
- |
  unswathe
- |
  unswayed
- |
  unsweetened
- |
  unswerving
- |
  unswervingly
- |
  unsystematic
- |
  untactful
- |
  untactfully
- |
  untainted
- |
  untalented
- |
  untamed
- |
  untangle
- |
  untanned
- |
  untapped
- |
  untarnished
- |
  untasted
- |
  untasteful
- |
  untaught
- |
  untaxed
- |
  unteachable
- |
  untempted
- |
  untempting
- |
  untenable
- |
  untenanted
- |
  untended
- |
  untested
- |
  unthankful
- |
  unthinkable
- |
  unthinkably
- |
  unthinking
- |
  unthinkingly
- |
  unthought
- |
  unthoughtful
- |
  unthrifty
- |
  unthrone
- |
  untidily
- |
  untidiness
- |
  untidy
- |
  untie
- |
  until
- |
  untilled
- |
  untimeliness
- |
  untimely
- |
  untired
- |
  untiring
- |
  untiringly
- |
  untitled
- |
  untold
- |
  Untouchable
- |
  untouchable
- |
  untouched
- |
  untoward
- |
  untowardly
- |
  untowardness
- |
  untraceable
- |
  untractable
- |
  untrained
- |
  untrammeled
- |
  untrammelled
- |
  untranslated
- |
  untraveled
- |
  untravelled
- |
  untraversed
- |
  untreated
- |
  untried
- |
  untrimmed
- |
  untrod
- |
  untrodden
- |
  untroubled
- |
  untrue
- |
  untrustful
- |
  untruth
- |
  untruthful
- |
  untruthfully
- |
  untune
- |
  untutored
- |
  untwine
- |
  untwist
- |
  untypical
- |
  unusable
- |
  unused
- |
  unusual
- |
  unusually
- |
  unutilized
- |
  unutterable
- |
  unutterably
- |
  unuttered
- |
  unvaried
- |
  unvarnished
- |
  unvarying
- |
  unveil
- |
  unveiling
- |
  unventilated
- |
  unverifiable
- |
  unverified
- |
  unversed
- |
  unvisited
- |
  unvoiced
- |
  unwanted
- |
  unwarily
- |
  unwariness
- |
  unwarmed
- |
  unwarranted
- |
  unwary
- |
  unwashed
- |
  unwatched
- |
  unwavering
- |
  unwaveringly
- |
  unweaned
- |
  unwearable
- |
  unwearied
- |
  unwearying
- |
  unweathered
- |
  unweave
- |
  unwed
- |
  unwelcome
- |
  unwell
- |
  unwholesome
- |
  unwieldily
- |
  unwieldiness
- |
  unwieldy
- |
  unwilling
- |
  unwillingly
- |
  unwind
- |
  unwise
- |
  unwisely
- |
  unwitnessed
- |
  unwitting
- |
  unwittingly
- |
  unwomanly
- |
  unwon
- |
  unwonted
- |
  unwontedly
- |
  unworkable
- |
  unworkably
- |
  unworldly
- |
  unworn
- |
  unworried
- |
  unworthily
- |
  unworthiness
- |
  unworthy
- |
  unwound
- |
  unwounded
- |
  unwove
- |
  unwoven
- |
  unwrap
- |
  unwrinkled
- |
  unwritten
- |
  unyielding
- |
  unyoke
- |
  unzip
- |
  Upanishad
- |
  upbeat
- |
  upbraid
- |
  upbringing
- |
  upchuck
- |
  upcoming
- |
  upcountry
- |
  update
- |
  Updike
- |
  updraft
- |
  upend
- |
  upfront
- |
  upgrade
- |
  upgrowth
- |
  upheaval
- |
  upheld
- |
  uphill
- |
  uphold
- |
  upholder
- |
  upholster
- |
  upholstered
- |
  upholsterer
- |
  upholstery
- |
  upkeep
- |
  upland
- |
  uplift
- |
  uplifting
- |
  upload
- |
  upmarket
- |
  upmost
- |
  Upper
- |
  upper
- |
  uppercase
- |
  uppercut
- |
  uppermost
- |
  uppish
- |
  uppishly
- |
  uppishness
- |
  uppity
- |
  Uppsala
- |
  upraise
- |
  uprear
- |
  upright
- |
  uprightly
- |
  uprightness
- |
  uprising
- |
  upriver
- |
  uproar
- |
  uproarious
- |
  uproariously
- |
  uproot
- |
  uprootedness
- |
  upscale
- |
  upset
- |
  upsetting
- |
  upshot
- |
  upside
- |
  upsilon
- |
  upstage
- |
  upstairs
- |
  upstanding
- |
  upstart
- |
  upstate
- |
  upstream
- |
  upstroke
- |
  upsurge
- |
  upsweep
- |
  upswept
- |
  upswing
- |
  uptake
- |
  uptalk
- |
  uptempo
- |
  upthrust
- |
  uptick
- |
  uptight
- |
  uptown
- |
  upturn
- |
  upturned
- |
  upward
- |
  upwardly
- |
  upwards
- |
  upwell
- |
  upwelling
- |
  upwind
- |
  uracil
- |
  Uralian
- |
  Uralic
- |
  Urals
- |
  uranium
- |
  uranographer
- |
  uranographic
- |
  uranography
- |
  Uranus
- |
  Urban
- |
  urban
- |
  urbane
- |
  urbanely
- |
  urbanisation
- |
  urbanite
- |
  urbanity
- |
  urbanization
- |
  urbanize
- |
  urbanologist
- |
  urbanology
- |
  urchin
- |
  uremia
- |
  uremic
- |
  ureter
- |
  urethane
- |
  urethra
- |
  urethrae
- |
  urethral
- |
  urethritis
- |
  urgency
- |
  urgent
- |
  urgently
- |
  Uriah
- |
  Uriel
- |
  urinal
- |
  urinalyses
- |
  urinalysis
- |
  urinary
- |
  urinate
- |
  urination
- |
  urine
- |
  urogenital
- |
  urologic
- |
  urological
- |
  urologist
- |
  urology
- |
  ursine
- |
  Ursula
- |
  urtext
- |
  urtexte
- |
  urticaria
- |
  urticate
- |
  urticating
- |
  urtication
- |
  Uruguay
- |
  Uruguayan
- |
  Urumchi
- |
  Urumqi
- |
  usability
- |
  usable
- |
  usably
- |
  usage
- |
  useability
- |
  useable
- |
  useful
- |
  usefully
- |
  usefulness
- |
  useless
- |
  uselessly
- |
  uselessness
- |
  USENET
- |
  Usenet
- |
  username
- |
  usher
- |
  usherette
- |
  Uspallata
- |
  Ustinov
- |
  usual
- |
  usually
- |
  usualness
- |
  usufruct
- |
  usurer
- |
  usurious
- |
  usuriously
- |
  usuriousness
- |
  usurp
- |
  usurpation
- |
  usurper
- |
  usury
- |
  Utahan
- |
  Utahn
- |
  utensil
- |
  uteri
- |
  uterine
- |
  uterus
- |
  utile
- |
  utilise
- |
  utilitarian
- |
  utilities
- |
  utility
- |
  utilizable
- |
  utilization
- |
  utilize
- |
  utilizer
- |
  utmost
- |
  Utopia
- |
  utopia
- |
  Utopian
- |
  utopian
- |
  Utrecht
- |
  Utrillo
- |
  utter
- |
  utterable
- |
  utterance
- |
  utterer
- |
  utterly
- |
  uttermost
- |
  uvula
- |
  uvulae
- |
  uvular
- |
  uxorial
- |
  uxorious
- |
  uxoriously
- |
  uxoriousness
- |
  Uzbek
- |
  Uzbekistan
- |
  vacancy
- |
  vacant
- |
  vacantly
- |
  vacate
- |
  vacation
- |
  vacationer
- |
  vacationist
- |
  vacationland
- |
  vaccinate
- |
  vaccination
- |
  vaccinator
- |
  vaccine
- |
  vaccinia
- |
  vacillate
- |
  vacillation
- |
  vacillator
- |
  vacua
- |
  vacuity
- |
  vacuolar
- |
  vacuole
- |
  vacuous
- |
  vacuously
- |
  vacuousness
- |
  vacuum
- |
  Vaduz
- |
  vagabond
- |
  vagabondage
- |
  vagaries
- |
  vagarious
- |
  vagariously
- |
  vagary
- |
  vagina
- |
  vaginae
- |
  vaginal
- |
  vaginitis
- |
  vagrancy
- |
  vagrant
- |
  vagrantly
- |
  vague
- |
  vaguely
- |
  vagueness
- |
  vainglorious
- |
  vainglory
- |
  vainly
- |
  valance
- |
  valanced
- |
  Valdez
- |
  valediction
- |
  valedictory
- |
  valence
- |
  Valencia
- |
  Valenciennes
- |
  valency
- |
  Valentine
- |
  valentine
- |
  Valentino
- |
  Valerian
- |
  valerian
- |
  Valerie
- |
  Valery
- |
  valet
- |
  Valhalla
- |
  valiance
- |
  valiant
- |
  valiantly
- |
  valid
- |
  validate
- |
  validation
- |
  validity
- |
  validly
- |
  validness
- |
  valise
- |
  Valium
- |
  Valkyrie
- |
  Valladolid
- |
  Vallejo
- |
  Valletta
- |
  valley
- |
  valor
- |
  valorization
- |
  valorize
- |
  valorous
- |
  valour
- |
  Valparaiso
- |
  valse
- |
  valuable
- |
  valuables
- |
  valuably
- |
  valuate
- |
  valuation
- |
  valuator
- |
  value
- |
  valued
- |
  valueless
- |
  valuer
- |
  values
- |
  valve
- |
  valved
- |
  valveless
- |
  valvular
- |
  vamoose
- |
  vamper
- |
  vampire
- |
  vampish
- |
  vampishly
- |
  vampy
- |
  vanadium
- |
  Vance
- |
  Vancouver
- |
  Vandal
- |
  vandal
- |
  vandalise
- |
  vandalism
- |
  vandalize
- |
  Vanderbilt
- |
  Vandyke
- |
  Vanessa
- |
  vanguard
- |
  vanguardism
- |
  vanguardist
- |
  vanilla
- |
  vanillin
- |
  vanish
- |
  vanisher
- |
  vanishing
- |
  vanity
- |
  vanquish
- |
  vanquisher
- |
  vantage
- |
  Vanuatu
- |
  Vanuatuan
- |
  Vanzetti
- |
  vapid
- |
  vapidity
- |
  vapidly
- |
  vapidness
- |
  vapor
- |
  vaporing
- |
  vaporise
- |
  vaporization
- |
  vaporize
- |
  vaporizer
- |
  vaporous
- |
  vaporously
- |
  vaporousness
- |
  vapors
- |
  vaporware
- |
  vapory
- |
  vapour
- |
  vaquero
- |
  Varanasi
- |
  variability
- |
  variable
- |
  variableness
- |
  variables
- |
  variably
- |
  variance
- |
  variant
- |
  variation
- |
  varicolored
- |
  varicose
- |
  varicosed
- |
  varicosity
- |
  varied
- |
  variedly
- |
  variegate
- |
  variegated
- |
  variegation
- |
  varietal
- |
  varietally
- |
  variety
- |
  variorum
- |
  various
- |
  variously
- |
  varlet
- |
  varletry
- |
  varment
- |
  varmint
- |
  Varna
- |
  varnish
- |
  varsity
- |
  varying
- |
  Vasari
- |
  vascular
- |
  vascularity
- |
  vasectomize
- |
  vasectomy
- |
  Vaseline
- |
  vasodilation
- |
  vasodilator
- |
  vasomotor
- |
  vassal
- |
  vassalage
- |
  vastly
- |
  vastness
- |
  vasty
- |
  vatic
- |
  Vatican
- |
  vaticinal
- |
  vaticinate
- |
  vaticination
- |
  vaticinator
- |
  vaticinatory
- |
  vaudeville
- |
  vaudevillian
- |
  Vaughan
- |
  Vaughn
- |
  vault
- |
  vaulted
- |
  vaulter
- |
  vaulting
- |
  vaulty
- |
  vaunt
- |
  vaunted
- |
  vaunter
- |
  vauntingly
- |
  Veadar
- |
  Veblen
- |
  vector
- |
  Vedanta
- |
  Vedantic
- |
  vedette
- |
  Vedic
- |
  vedic
- |
  veejay
- |
  vegan
- |
  veganism
- |
  vegetable
- |
  vegetal
- |
  vegetarian
- |
  vegetate
- |
  vegetation
- |
  vegetational
- |
  vegetative
- |
  vegetatively
- |
  veggie
- |
  veggies
- |
  vehemence
- |
  vehemency
- |
  vehement
- |
  vehemently
- |
  vehicle
- |
  vehicular
- |
  veiled
- |
  veined
- |
  veining
- |
  veiny
- |
  velar
- |
  Velazquez
- |
  Velcro
- |
  veldt
- |
  velleity
- |
  vellum
- |
  Velma
- |
  velocipede
- |
  velocity
- |
  velodrome
- |
  velour
- |
  velours
- |
  velum
- |
  velutinous
- |
  velvet
- |
  velveteen
- |
  velvety
- |
  venal
- |
  venality
- |
  venally
- |
  venation
- |
  venational
- |
  vendee
- |
  vender
- |
  vendetta
- |
  vendible
- |
  vendor
- |
  veneer
- |
  veneered
- |
  venerability
- |
  venerable
- |
  venerably
- |
  venerate
- |
  venerated
- |
  veneration
- |
  venerator
- |
  venereal
- |
  venereally
- |
  venery
- |
  Venetian
- |
  Venezia
- |
  Venezuela
- |
  Venezuelan
- |
  vengeance
- |
  vengeful
- |
  vengefully
- |
  vengefulness
- |
  venial
- |
  veniality
- |
  venially
- |
  Venice
- |
  venire
- |
  venireman
- |
  venison
- |
  venom
- |
  venomous
- |
  venomously
- |
  venomousness
- |
  venosity
- |
  venous
- |
  venously
- |
  ventilate
- |
  ventilated
- |
  ventilation
- |
  ventilator
- |
  ventral
- |
  ventrally
- |
  ventricle
- |
  ventricular
- |
  ventriloquy
- |
  Ventura
- |
  venture
- |
  venturesome
- |
  venturous
- |
  venturously
- |
  venue
- |
  Venus
- |
  Venusian
- |
  veracious
- |
  veraciously
- |
  veracity
- |
  Veracruz
- |
  veranda
- |
  verandah
- |
  verbal
- |
  verbalism
- |
  verbalist
- |
  verbalistic
- |
  verbalizable
- |
  verbalize
- |
  verbalizer
- |
  verbally
- |
  verbatim
- |
  verbena
- |
  verbiage
- |
  verbose
- |
  verbosely
- |
  verbosity
- |
  verboten
- |
  verdancy
- |
  verdant
- |
  verdantly
- |
  Verde
- |
  Verdi
- |
  verdict
- |
  verdigris
- |
  Verdun
- |
  verdure
- |
  verdured
- |
  verdurous
- |
  verge
- |
  verger
- |
  Vergil
- |
  veridical
- |
  veridicality
- |
  veridically
- |
  verifiable
- |
  verifiably
- |
  verification
- |
  verifier
- |
  verify
- |
  verily
- |
  verisimilar
- |
  verism
- |
  verismo
- |
  verist
- |
  veristic
- |
  veritable
- |
  veritably
- |
  verite
- |
  verity
- |
  Vermeer
- |
  vermeil
- |
  vermicelli
- |
  vermicide
- |
  vermiculite
- |
  vermiform
- |
  vermifuge
- |
  vermilion
- |
  vermillion
- |
  vermin
- |
  verminous
- |
  Vermont
- |
  Vermonter
- |
  vermouth
- |
  Verna
- |
  vernacular
- |
  vernacularly
- |
  vernal
- |
  vernally
- |
  Verne
- |
  vernier
- |
  Vernon
- |
  Verona
- |
  Veronese
- |
  Veronica
- |
  veronica
- |
  Verrazano
- |
  Verrazzano
- |
  Versailles
- |
  versatile
- |
  versatilely
- |
  versatility
- |
  verse
- |
  versed
- |
  versicle
- |
  versifier
- |
  versify
- |
  version
- |
  verso
- |
  versus
- |
  vertebra
- |
  vertebrae
- |
  vertebral
- |
  vertebrate
- |
  vertex
- |
  vertical
- |
  verticality
- |
  vertically
- |
  vertices
- |
  vertiginous
- |
  vertigo
- |
  vertu
- |
  vervain
- |
  verve
- |
  vesicant
- |
  vesicle
- |
  vesicular
- |
  vesiculate
- |
  vesiculated
- |
  vesiculation
- |
  Vespasian
- |
  vesper
- |
  Vespers
- |
  vespers
- |
  vespertine
- |
  vespine
- |
  Vespucci
- |
  vessel
- |
  Vesta
- |
  vestal
- |
  vested
- |
  vestiary
- |
  vestibular
- |
  vestibule
- |
  vestibuled
- |
  vestige
- |
  vestigial
- |
  vestigially
- |
  vesting
- |
  vestment
- |
  vestments
- |
  vestry
- |
  vestryman
- |
  vesture
- |
  Vesuvian
- |
  Vesuvius
- |
  vetch
- |
  veteran
- |
  veterinarian
- |
  veterinary
- |
  vetoer
- |
  vetting
- |
  vexation
- |
  vexatious
- |
  vexatiously
- |
  vexed
- |
  vexillology
- |
  viability
- |
  viable
- |
  viably
- |
  viaduct
- |
  viand
- |
  viands
- |
  viatica
- |
  viaticum
- |
  vibes
- |
  vibraharp
- |
  vibrancy
- |
  vibrant
- |
  vibrantly
- |
  vibraphone
- |
  vibraphonist
- |
  vibrate
- |
  vibration
- |
  vibrational
- |
  vibrations
- |
  vibrato
- |
  vibrator
- |
  vibratory
- |
  viburnum
- |
  vicar
- |
  vicarage
- |
  vicariate
- |
  vicarious
- |
  vicariously
- |
  vicarship
- |
  vicegerency
- |
  vicegerent
- |
  vicennial
- |
  viceregal
- |
  viceroy
- |
  viceroyal
- |
  viceroyalty
- |
  viceroyship
- |
  Vichy
- |
  vichyssoise
- |
  vicinage
- |
  vicinal
- |
  vicinity
- |
  vicious
- |
  viciously
- |
  viciousness
- |
  vicissitude
- |
  vicissitudes
- |
  Vicki
- |
  Vickie
- |
  Vicksburg
- |
  Vicky
- |
  victim
- |
  victimise
- |
  victimize
- |
  victimizer
- |
  victimless
- |
  Victor
- |
  victor
- |
  Victoria
- |
  victoria
- |
  Victorian
- |
  Victorianism
- |
  victorious
- |
  victoriously
- |
  victory
- |
  victual
- |
  victualer
- |
  victualler
- |
  victuals
- |
  vicuna
- |
  Vidal
- |
  videlicet
- |
  video
- |
  videodisc
- |
  videodisk
- |
  videophone
- |
  videotape
- |
  Vienna
- |
  Viennese
- |
  Vientiane
- |
  Vietcong
- |
  Vietnam
- |
  Vietnamese
- |
  viewer
- |
  viewership
- |
  viewfinder
- |
  viewpoint
- |
  vigesimal
- |
  vigil
- |
  vigilance
- |
  vigilant
- |
  vigilante
- |
  vigilanteism
- |
  vigilantism
- |
  vigilantist
- |
  vigilantly
- |
  vigils
- |
  vignette
- |
  vignettist
- |
  vigor
- |
  vigorless
- |
  vigorous
- |
  vigorously
- |
  vigorousness
- |
  vigour
- |
  Vijayawada
- |
  Viking
- |
  viking
- |
  vilely
- |
  vileness
- |
  vilification
- |
  vilifier
- |
  vilify
- |
  Villa
- |
  villa
- |
  village
- |
  villager
- |
  Villahermosa
- |
  villain
- |
  villainess
- |
  villainous
- |
  villainously
- |
  villainy
- |
  villein
- |
  villeinage
- |
  villi
- |
  Villon
- |
  villous
- |
  villus
- |
  Vilna
- |
  Vilnius
- |
  vinaigrette
- |
  Vincent
- |
  Vinci
- |
  vincible
- |
  vindicable
- |
  vindicate
- |
  vindication
- |
  vindicator
- |
  vindicatory
- |
  vindictive
- |
  vindictively
- |
  Vindobna
- |
  Vindobona
- |
  vinegar
- |
  vinegary
- |
  vineyard
- |
  vinicultural
- |
  viniculture
- |
  Vinland
- |
  vinosity
- |
  vinous
- |
  vinously
- |
  vintage
- |
  vintner
- |
  vinyl
- |
  Viola
- |
  viola
- |
  violable
- |
  violate
- |
  violation
- |
  violative
- |
  violator
- |
  violence
- |
  violent
- |
  violently
- |
  Violet
- |
  violet
- |
  violin
- |
  violinist
- |
  violist
- |
  violoncello
- |
  viper
- |
  viperine
- |
  viperish
- |
  viperous
- |
  virago
- |
  viral
- |
  virally
- |
  vireo
- |
  virescence
- |
  virescent
- |
  virescently
- |
  Virgil
- |
  Virgilian
- |
  Virgin
- |
  virgin
- |
  virginal
- |
  virginally
- |
  Virginia
- |
  Virginian
- |
  virginity
- |
  Virgo
- |
  virgule
- |
  viridescence
- |
  viridescent
- |
  viridity
- |
  virile
- |
  virility
- |
  virion
- |
  virologist
- |
  virology
- |
  virtu
- |
  virtual
- |
  virtuality
- |
  virtually
- |
  virtue
- |
  virtueless
- |
  virtues
- |
  virtuosi
- |
  virtuosic
- |
  virtuosity
- |
  virtuoso
- |
  virtuous
- |
  virtuously
- |
  virtuousness
- |
  virulence
- |
  virulent
- |
  virulently
- |
  virus
- |
  visage
- |
  visaged
- |
  Visayan
- |
  viscera
- |
  visceral
- |
  viscerally
- |
  viscid
- |
  viscidity
- |
  viscidly
- |
  viscose
- |
  viscosity
- |
  viscount
- |
  viscountcy
- |
  viscountess
- |
  viscous
- |
  viscously
- |
  viscousness
- |
  viscus
- |
  Vishnu
- |
  visibility
- |
  visible
- |
  visibly
- |
  Visigoth
- |
  vision
- |
  visionary
- |
  visit
- |
  visitable
- |
  visitant
- |
  visitation
- |
  visitational
- |
  visitor
- |
  visor
- |
  visored
- |
  vista
- |
  Vistula
- |
  visual
- |
  visualise
- |
  visualize
- |
  visualizer
- |
  visually
- |
  vitae
- |
  vital
- |
  vitalism
- |
  vitalist
- |
  vitalistic
- |
  vitality
- |
  vitalization
- |
  vitalize
- |
  vitalizer
- |
  vitally
- |
  vitals
- |
  vitamin
- |
  vitiate
- |
  vitiation
- |
  vitiator
- |
  viticultural
- |
  viticulture
- |
  vitreous
- |
  vitreousness
- |
  vitrifaction
- |
  vitrifiable
- |
  vitrify
- |
  vitrine
- |
  vitriol
- |
  vitriolic
- |
  Vitsyebsk
- |
  vittles
- |
  vituperate
- |
  vituperation
- |
  vituperative
- |
  vituperator
- |
  vivace
- |
  vivacious
- |
  vivaciously
- |
  vivacity
- |
  Vivaldi
- |
  Vivian
- |
  vivid
- |
  vividly
- |
  vividness
- |
  vivification
- |
  vivifier
- |
  vivify
- |
  viviparity
- |
  viviparous
- |
  viviparously
- |
  vivisect
- |
  vivisection
- |
  vivisector
- |
  vixen
- |
  vixenish
- |
  vixenishly
- |
  vizard
- |
  vizier
- |
  vizierate
- |
  vizierial
- |
  viziership
- |
  vizir
- |
  vizor
- |
  Vladikavkaz
- |
  Vladivostok
- |
  Vlaminck
- |
  vocable
- |
  vocabulary
- |
  vocal
- |
  vocalic
- |
  vocalist
- |
  vocalization
- |
  vocalize
- |
  vocalizer
- |
  vocally
- |
  vocals
- |
  vocation
- |
  vocational
- |
  vocationally
- |
  vocative
- |
  vociferant
- |
  vociferate
- |
  vociferation
- |
  vociferator
- |
  vociferous
- |
  vociferously
- |
  vodka
- |
  vogue
- |
  voguish
- |
  voice
- |
  voiced
- |
  voicedness
- |
  voiceless
- |
  voicelessly
- |
  voiceover
- |
  voiceprint
- |
  voidable
- |
  voider
- |
  voila
- |
  voile
- |
  Volans
- |
  volant
- |
  volatile
- |
  volatiles
- |
  volatility
- |
  volatilize
- |
  volcanic
- |
  volcanically
- |
  volcanism
- |
  volcano
- |
  volcanology
- |
  Volga
- |
  Volgograd
- |
  volitant
- |
  volition
- |
  volitional
- |
  volitionally
- |
  volitive
- |
  volley
- |
  volleyball
- |
  volleyer
- |
  Volos
- |
  Volstead
- |
  Volta
- |
  voltage
- |
  voltaic
- |
  Voltaire
- |
  voltmeter
- |
  volubility
- |
  voluble
- |
  volubleness
- |
  volubly
- |
  volume
- |
  volumetric
- |
  voluminous
- |
  voluminously
- |
  voluntarily
- |
  voluntarism
- |
  voluntarist
- |
  voluntary
- |
  volunteer
- |
  volunteerism
- |
  voluptuary
- |
  voluptuous
- |
  voluptuously
- |
  volute
- |
  voluted
- |
  volution
- |
  vomit
- |
  vomiting
- |
  vomitous
- |
  Vonnegut
- |
  voodoo
- |
  voodooism
- |
  voracious
- |
  voraciously
- |
  voracity
- |
  Voronezh
- |
  vortex
- |
  vortical
- |
  vortically
- |
  vortices
- |
  vorticity
- |
  vorticose
- |
  vorticular
- |
  Vosges
- |
  votarist
- |
  votary
- |
  voteless
- |
  voter
- |
  voting
- |
  votive
- |
  vouch
- |
  voucher
- |
  vouchsafe
- |
  voussoir
- |
  vowel
- |
  vower
- |
  voyage
- |
  voyager
- |
  voyageur
- |
  voyaging
- |
  voyeur
- |
  voyeurism
- |
  voyeuristic
- |
  Vulcan
- |
  vulcanism
- |
  vulcanizable
- |
  vulcanize
- |
  vulcanizer
- |
  vulcanology
- |
  vulgar
- |
  vulgarian
- |
  vulgarism
- |
  vulgarity
- |
  vulgarize
- |
  vulgarizer
- |
  vulgarly
- |
  Vulgate
- |
  vulgate
- |
  vulnerable
- |
  vulnerably
- |
  Vulpecula
- |
  vulpine
- |
  vulture
- |
  vulturous
- |
  vulva
- |
  vulvae
- |
  vulval
- |
  vulvar
- |
  vying
- |
  Wabash
- |
  wabble
- |
  wackily
- |
  wackiness
- |
  wacko
- |
  wacky
- |
  wadable
- |
  wadding
- |
  waddle
- |
  waddler
- |
  wadeable
- |
  wader
- |
  waders
- |
  wafer
- |
  waffle
- |
  waffler
- |
  waffling
- |
  wager
- |
  wagerer
- |
  wages
- |
  waggery
- |
  waggish
- |
  waggishly
- |
  waggishness
- |
  waggle
- |
  waggly
- |
  waggon
- |
  Wagner
- |
  Wagnerian
- |
  wagon
- |
  wagoner
- |
  wagonette
- |
  wagtail
- |
  wahine
- |
  wahoo
- |
  waifish
- |
  Waikiki
- |
  wailer
- |
  wailful
- |
  wailfully
- |
  wailing
- |
  wainscot
- |
  wainscoting
- |
  wainscotting
- |
  wainwright
- |
  waist
- |
  waistband
- |
  waistcoat
- |
  waisted
- |
  waistline
- |
  waiter
- |
  waiting
- |
  waitperson
- |
  waitress
- |
  waitressing
- |
  waitron
- |
  waitstaff
- |
  waive
- |
  waiver
- |
  Wakefield
- |
  wakeful
- |
  wakefully
- |
  wakefulness
- |
  waken
- |
  wakener
- |
  waking
- |
  Walachia
- |
  Walcott
- |
  Waldheim
- |
  Waldo
- |
  Wales
- |
  Walesa
- |
  walkable
- |
  walkaway
- |
  Walker
- |
  walker
- |
  walking
- |
  walkingstick
- |
  Walkman
- |
  walkout
- |
  walkover
- |
  walkup
- |
  walkway
- |
  wallaby
- |
  Wallace
- |
  Wallachia
- |
  wallboard
- |
  walled
- |
  wallet
- |
  walleye
- |
  walleyed
- |
  wallflower
- |
  Wallis
- |
  Walloon
- |
  wallop
- |
  walloper
- |
  walloping
- |
  wallow
- |
  wallower
- |
  wallpaper
- |
  walls
- |
  walnut
- |
  Walpole
- |
  walrus
- |
  Walsall
- |
  Walter
- |
  Walton
- |
  waltz
- |
  waltzer
- |
  wamble
- |
  Wampanoag
- |
  wampum
- |
  Wanda
- |
  wander
- |
  wanderer
- |
  wanderingly
- |
  wanderlust
- |
  Wandsworth
- |
  wangle
- |
  wangler
- |
  Wankel
- |
  wanly
- |
  wanna
- |
  wannabe
- |
  wanness
- |
  wantad
- |
  wanted
- |
  wanting
- |
  wanton
- |
  wantonly
- |
  wantonness
- |
  wapiti
- |
  warble
- |
  warbler
- |
  warbonnet
- |
  warden
- |
  warder
- |
  wardrobe
- |
  wardroom
- |
  wardship
- |
  warehouse
- |
  warehouseman
- |
  warehouser
- |
  wareroom
- |
  wares
- |
  warfare
- |
  warfarin
- |
  warhead
- |
  Warhol
- |
  warhorse
- |
  warily
- |
  wariness
- |
  warless
- |
  Warley
- |
  warlike
- |
  warlock
- |
  warlord
- |
  warmblooded
- |
  warmer
- |
  warmhearted
- |
  warmish
- |
  warmly
- |
  warmness
- |
  warmonger
- |
  warmongering
- |
  warmth
- |
  Warner
- |
  warning
- |
  warningly
- |
  warpage
- |
  warpath
- |
  warped
- |
  warper
- |
  warplane
- |
  warrant
- |
  warrantable
- |
  warranted
- |
  warrantee
- |
  warranter
- |
  warranty
- |
  Warren
- |
  warren
- |
  warring
- |
  warrior
- |
  Warsaw
- |
  warship
- |
  warthog
- |
  wartime
- |
  warty
- |
  Warwick
- |
  Warwickshire
- |
  wasabi
- |
  Wasatch
- |
  washable
- |
  washbasin
- |
  washboard
- |
  washbowl
- |
  washcloth
- |
  washer
- |
  washerwoman
- |
  washhouse
- |
  washily
- |
  washiness
- |
  washing
- |
  Washington
- |
  washout
- |
  washrag
- |
  washroom
- |
  washstand
- |
  washtub
- |
  washwoman
- |
  washy
- |
  Waspish
- |
  waspish
- |
  waspishly
- |
  waspishness
- |
  Waspy
- |
  wassail
- |
  wassailer
- |
  wastage
- |
  waste
- |
  wastebasket
- |
  wasted
- |
  wasteful
- |
  wastefully
- |
  wastefulness
- |
  wasteland
- |
  wastepaper
- |
  waster
- |
  wastes
- |
  wastrel
- |
  watch
- |
  watchband
- |
  watchdog
- |
  watcher
- |
  watchful
- |
  watchfully
- |
  watchfulness
- |
  watchmaker
- |
  watchmaking
- |
  watchman
- |
  watchtower
- |
  watchword
- |
  water
- |
  waterbed
- |
  waterborne
- |
  Waterbury
- |
  watercolor
- |
  watercolour
- |
  watercourse
- |
  watercraft
- |
  watercress
- |
  waterfall
- |
  waterfowl
- |
  waterfront
- |
  Watergate
- |
  waterglass
- |
  waterhole
- |
  wateriness
- |
  waterish
- |
  waterlily
- |
  waterline
- |
  waterlogged
- |
  Waterloo
- |
  waterloo
- |
  waterman
- |
  watermark
- |
  watermelon
- |
  waterpower
- |
  waterproof
- |
  waters
- |
  watershed
- |
  waterside
- |
  waterspout
- |
  watertight
- |
  waterway
- |
  waterwheel
- |
  waterworks
- |
  watery
- |
  Watson
- |
  wattage
- |
  Watteau
- |
  wattle
- |
  wattled
- |
  wattles
- |
  Waugh
- |
  waveband
- |
  waveform
- |
  wavelength
- |
  wavelet
- |
  wavelike
- |
  waver
- |
  waverer
- |
  waveringly
- |
  Waverley
- |
  wavily
- |
  waviness
- |
  waxen
- |
  waxiness
- |
  waxwing
- |
  waxwork
- |
  waxworks
- |
  waybill
- |
  wayfarer
- |
  wayfaring
- |
  waylaid
- |
  waylay
- |
  waylayer
- |
  Wayne
- |
  wayside
- |
  wayward
- |
  waywardly
- |
  waywardness
- |
  weaken
- |
  weakener
- |
  weakfish
- |
  weakish
- |
  weakling
- |
  weakly
- |
  weakness
- |
  weald
- |
  wealth
- |
  wealthiness
- |
  wealthy
- |
  weaning
- |
  weapon
- |
  weaponless
- |
  weaponry
- |
  wearable
- |
  wearer
- |
  weariless
- |
  wearily
- |
  weariness
- |
  wearisome
- |
  wearisomely
- |
  weary
- |
  weasel
- |
  weaselly
- |
  weather
- |
  weatherboard
- |
  weathercock
- |
  weathered
- |
  weathering
- |
  weatherize
- |
  weatherman
- |
  weatherproof
- |
  weatherstrip
- |
  weathervane
- |
  weatherworn
- |
  weave
- |
  weaver
- |
  webbed
- |
  webbing
- |
  webcast
- |
  Weber
- |
  weber
- |
  webfeet
- |
  webfoot
- |
  webmaster
- |
  webpage
- |
  website
- |
  Webster
- |
  webworm
- |
  wedded
- |
  wedding
- |
  wedge
- |
  wedgie
- |
  Wedgwood
- |
  wedlock
- |
  Wednesday
- |
  weeder
- |
  weediness
- |
  weeding
- |
  weedless
- |
  weeds
- |
  weedy
- |
  weekday
- |
  weekend
- |
  weekly
- |
  weeknight
- |
  weenie
- |
  weensy
- |
  weeny
- |
  weeper
- |
  weeping
- |
  weepy
- |
  weevil
- |
  weevilly
- |
  weevily
- |
  weigh
- |
  weight
- |
  weighted
- |
  weightily
- |
  weightiness
- |
  weightless
- |
  weightlessly
- |
  weightlifter
- |
  weighty
- |
  Weill
- |
  Weimar
- |
  weird
- |
  weirdie
- |
  weirdly
- |
  weirdness
- |
  weirdo
- |
  Weizmann
- |
  Welch
- |
  welch
- |
  welcome
- |
  weldable
- |
  welder
- |
  welding
- |
  Weldon
- |
  Welfare
- |
  welfare
- |
  welkin
- |
  Welland
- |
  wellborn
- |
  Welles
- |
  wellhead
- |
  Wellington
- |
  wellness
- |
  Wells
- |
  wellspring
- |
  Welsh
- |
  welsh
- |
  welsher
- |
  Welshman
- |
  Welshwoman
- |
  welter
- |
  welterweight
- |
  Welty
- |
  wench
- |
  Wendell
- |
  wendigo
- |
  Wendy
- |
  werewolf
- |
  werewolves
- |
  Werner
- |
  werwolf
- |
  Weser
- |
  weskit
- |
  Wesley
- |
  Wesleyan
- |
  Wessex
- |
  westbound
- |
  westerlies
- |
  westerly
- |
  Western
- |
  western
- |
  Westerner
- |
  westerner
- |
  westernize
- |
  westernmost
- |
  Westinghouse
- |
  Westminster
- |
  Westphalia
- |
  Westphalian
- |
  westward
- |
  westwardly
- |
  westwards
- |
  wetback
- |
  wether
- |
  wetland
- |
  wetlands
- |
  wetly
- |
  wetness
- |
  wetsuit
- |
  wetter
- |
  Weyden
- |
  whack
- |
  whacked
- |
  whacker
- |
  whacky
- |
  whale
- |
  whaleboat
- |
  whalebone
- |
  whaler
- |
  whaling
- |
  whammy
- |
  wharf
- |
  wharfage
- |
  Wharton
- |
  wharves
- |
  whatever
- |
  whatnot
- |
  whatsoever
- |
  wheal
- |
  wheat
- |
  wheaten
- |
  Wheatley
- |
  Wheatstone
- |
  wheedle
- |
  wheedler
- |
  wheedlingly
- |
  wheel
- |
  wheelbarrow
- |
  wheelbase
- |
  wheelchair
- |
  wheeled
- |
  wheeler
- |
  wheelhorse
- |
  wheelhouse
- |
  wheelie
- |
  Wheeling
- |
  wheelless
- |
  wheels
- |
  wheelwright
- |
  wheeze
- |
  wheezer
- |
  wheezily
- |
  wheeziness
- |
  wheezy
- |
  whelk
- |
  whelm
- |
  whelp
- |
  whence
- |
  whenever
- |
  whensoever
- |
  where
- |
  whereabout
- |
  whereabouts
- |
  whereas
- |
  whereat
- |
  whereby
- |
  wherefore
- |
  wherein
- |
  whereof
- |
  whereon
- |
  wheresoever
- |
  whereto
- |
  whereupon
- |
  wherever
- |
  wherewith
- |
  wherewithal
- |
  wherry
- |
  wherryman
- |
  whether
- |
  whetstone
- |
  whetter
- |
  which
- |
  whichever
- |
  whichsoever
- |
  whicker
- |
  whiff
- |
  whiffletree
- |
  Whiggery
- |
  Whiggish
- |
  Whiggism
- |
  while
- |
  whilom
- |
  whilst
- |
  whimper
- |
  whimperingly
- |
  whimsey
- |
  whimsical
- |
  whimsicality
- |
  whimsically
- |
  whimsy
- |
  whine
- |
  whiner
- |
  whiney
- |
  whinge
- |
  whingeingly
- |
  whinger
- |
  whingy
- |
  whinny
- |
  whiny
- |
  whipcord
- |
  whiplash
- |
  whipper
- |
  whippet
- |
  whipping
- |
  whippletree
- |
  whippoorwill
- |
  whipsaw
- |
  whipstitch
- |
  whipt
- |
  whirl
- |
  whirler
- |
  whirligig
- |
  whirlpool
- |
  whirlwind
- |
  whirlybird
- |
  whirr
- |
  whish
- |
  whisk
- |
  whiskbroom
- |
  whisker
- |
  whiskered
- |
  whiskers
- |
  whiskery
- |
  whiskey
- |
  whisky
- |
  whisper
- |
  whispered
- |
  whisperer
- |
  whispering
- |
  whispery
- |
  whist
- |
  whistle
- |
  Whistler
- |
  whistler
- |
  whistling
- |
  White
- |
  white
- |
  whitebait
- |
  whitecap
- |
  whitefish
- |
  Whitehall
- |
  Whitehead
- |
  whitehead
- |
  Whitehorse
- |
  whiten
- |
  whitener
- |
  whiteness
- |
  whitening
- |
  whiteout
- |
  whitepine
- |
  whites
- |
  whitetail
- |
  whitewall
- |
  whitewash
- |
  whitewasher
- |
  whitewater
- |
  whitewood
- |
  whither
- |
  whiting
- |
  whitish
- |
  whitlow
- |
  Whitman
- |
  Whitney
- |
  Whitsunday
- |
  Whittier
- |
  whittle
- |
  whittler
- |
  whizz
- |
  whodunit
- |
  whodunnit
- |
  whoever
- |
  whole
- |
  wholehearted
- |
  wholemeal
- |
  wholeness
- |
  wholesale
- |
  wholesaler
- |
  wholesome
- |
  wholesomely
- |
  wholism
- |
  wholistic
- |
  wholly
- |
  whomever
- |
  whomsoever
- |
  whoop
- |
  whooper
- |
  whoopla
- |
  whoops
- |
  whoosh
- |
  whopper
- |
  whopping
- |
  whore
- |
  whoreish
- |
  whorish
- |
  whorl
- |
  whorled
- |
  whose
- |
  whosesoever
- |
  whosever
- |
  whoso
- |
  whosoever
- |
  Wicca
- |
  Wiccan
- |
  Wichita
- |
  wicked
- |
  wickedly
- |
  wickedness
- |
  wicker
- |
  wickerwork
- |
  wicket
- |
  wickiup
- |
  widdershins
- |
  widely
- |
  widemouthed
- |
  widen
- |
  widener
- |
  wideness
- |
  widening
- |
  widespread
- |
  widgeon
- |
  widget
- |
  widow
- |
  widowed
- |
  widower
- |
  widowhood
- |
  width
- |
  widthways
- |
  widthwise
- |
  wield
- |
  wielder
- |
  wieldy
- |
  wiener
- |
  wienie
- |
  Wiesbaden
- |
  Wiesel
- |
  wifehood
- |
  wifeless
- |
  wifely
- |
  wigeon
- |
  wiggle
- |
  wiggler
- |
  wiggly
- |
  Wight
- |
  wight
- |
  wiglet
- |
  wigwag
- |
  wigwam
- |
  Wilber
- |
  Wilberforce
- |
  Wilbert
- |
  Wilbur
- |
  Wilda
- |
  wildcat
- |
  wildcatter
- |
  Wilde
- |
  wildebeest
- |
  Wilder
- |
  wilderness
- |
  wildfire
- |
  wildflower
- |
  wildfowl
- |
  wilding
- |
  wildlife
- |
  wildling
- |
  wildly
- |
  wildness
- |
  wilds
- |
  wildwood
- |
  wiles
- |
  Wiley
- |
  Wilford
- |
  Wilfred
- |
  wilful
- |
  wilfully
- |
  wilfulness
- |
  Wilhelm
- |
  Wilhelmina
- |
  wilily
- |
  wiliness
- |
  Wilkins
- |
  Willa
- |
  Willard
- |
  willed
- |
  Willemstad
- |
  willful
- |
  willfully
- |
  willfulness
- |
  William
- |
  Williams
- |
  Williamsburg
- |
  Willie
- |
  willies
- |
  willing
- |
  willingly
- |
  willingness
- |
  Willis
- |
  williwaw
- |
  willow
- |
  willowware
- |
  willowy
- |
  willpower
- |
  willywaw
- |
  Wilma
- |
  Wilmer
- |
  Wilmington
- |
  Wilson
- |
  Wilsonian
- |
  Wilton
- |
  Wiltshire
- |
  wimble
- |
  wimpish
- |
  wimpishly
- |
  wimpishness
- |
  wimple
- |
  wimpled
- |
  wimpy
- |
  wince
- |
  winch
- |
  Winchester
- |
  windage
- |
  windbag
- |
  windblown
- |
  windbreak
- |
  windbreaker
- |
  windburn
- |
  windburned
- |
  windchill
- |
  winded
- |
  winder
- |
  Windermere
- |
  windfall
- |
  windflower
- |
  Windhoek
- |
  windigo
- |
  windily
- |
  windiness
- |
  winding
- |
  windjammer
- |
  windlass
- |
  windless
- |
  windmill
- |
  window
- |
  windowdress
- |
  windowless
- |
  windowpane
- |
  Windows
- |
  windowsill
- |
  windpipe
- |
  windproof
- |
  windrow
- |
  winds
- |
  windscreen
- |
  windshield
- |
  windsock
- |
  Windsor
- |
  windstorm
- |
  windsurf
- |
  windsurfer
- |
  windsurfing
- |
  windswept
- |
  windup
- |
  windward
- |
  windy
- |
  wineglass
- |
  winegrower
- |
  winepress
- |
  winery
- |
  wineskin
- |
  Winfield
- |
  Winfred
- |
  wingding
- |
  winged
- |
  winger
- |
  wingless
- |
  winglike
- |
  wings
- |
  wingspan
- |
  wingspread
- |
  wingtip
- |
  Winifred
- |
  winker
- |
  winnable
- |
  Winnebago
- |
  winner
- |
  Winnie
- |
  winning
- |
  winningly
- |
  winnings
- |
  Winnipeg
- |
  Winnipegger
- |
  winnow
- |
  winnower
- |
  winsome
- |
  winsomely
- |
  winsomeness
- |
  Winston
- |
  winter
- |
  wintergreen
- |
  winterize
- |
  winterkill
- |
  wintertide
- |
  wintertime
- |
  wintery
- |
  Winthrop
- |
  Winton
- |
  wintriness
- |
  wintry
- |
  wiper
- |
  wired
- |
  wirehair
- |
  wirehaired
- |
  wireless
- |
  Wirephoto
- |
  wiretap
- |
  wiretapper
- |
  wiretapping
- |
  wireworm
- |
  wiriness
- |
  wiring
- |
  Wisconsin
- |
  Wisconsinite
- |
  Wisdom
- |
  wisdom
- |
  wiseacre
- |
  wisecrack
- |
  wisely
- |
  wisenheimer
- |
  wishbone
- |
  wisher
- |
  wishful
- |
  wishfully
- |
  wishfulness
- |
  wispy
- |
  wistaria
- |
  wisteria
- |
  wistful
- |
  wistfully
- |
  wistfulness
- |
  witch
- |
  witchcraft
- |
  witchery
- |
  witchgrass
- |
  witching
- |
  witchy
- |
  withal
- |
  withdraw
- |
  withdrawal
- |
  withdrawn
- |
  withdrew
- |
  withe
- |
  wither
- |
  withered
- |
  withering
- |
  witheringly
- |
  withers
- |
  withershins
- |
  withheld
- |
  withhold
- |
  withholding
- |
  within
- |
  without
- |
  withstand
- |
  withstood
- |
  withy
- |
  witless
- |
  witlessly
- |
  witlessness
- |
  witness
- |
  witted
- |
  Wittgenstein
- |
  witticism
- |
  wittily
- |
  wittiness
- |
  witting
- |
  wittingly
- |
  witty
- |
  wives
- |
  wizard
- |
  wizardly
- |
  wizardry
- |
  wizen
- |
  wizened
- |
  wobble
- |
  wobbliness
- |
  wobbly
- |
  Wodehouse
- |
  Woden
- |
  woebegone
- |
  woeful
- |
  woefully
- |
  woefulness
- |
  woful
- |
  woken
- |
  Wolfe
- |
  wolfhound
- |
  wolfish
- |
  wolfishly
- |
  wolfram
- |
  Wollaston
- |
  Wollongong
- |
  Wolsey
- |
  wolverine
- |
  wolves
- |
  woman
- |
  womanhood
- |
  womanish
- |
  womanize
- |
  womanizer
- |
  womankind
- |
  womanlike
- |
  womanliness
- |
  womanly
- |
  wombat
- |
  women
- |
  womenfolk
- |
  womenfolks
- |
  womenkind
- |
  Wonder
- |
  wonder
- |
  wonderful
- |
  wonderfully
- |
  wonderland
- |
  wonderment
- |
  wondrous
- |
  wondrously
- |
  wondrousness
- |
  wonted
- |
  wonton
- |
  woodbine
- |
  woodblock
- |
  woodcarver
- |
  woodcarving
- |
  woodchopper
- |
  woodchuck
- |
  woodcock
- |
  woodcraft
- |
  woodcut
- |
  woodcutter
- |
  woodcutting
- |
  wooded
- |
  wooden
- |
  woodenly
- |
  woodenness
- |
  woodenware
- |
  Woodhull
- |
  woodiness
- |
  woodland
- |
  woodlot
- |
  woodman
- |
  woodnote
- |
  woodpecker
- |
  woodpile
- |
  Woodrow
- |
  woodruff
- |
  Woods
- |
  woods
- |
  woodshed
- |
  woodsiness
- |
  woodsman
- |
  Woodstock
- |
  woodsy
- |
  woodwind
- |
  woodwork
- |
  woodworker
- |
  woodworking
- |
  woody
- |
  wooer
- |
  woofer
- |
  wooing
- |
  wooled
- |
  woolen
- |
  woolens
- |
  Woolf
- |
  woolgather
- |
  woolie
- |
  woollen
- |
  woolliness
- |
  woolly
- |
  wooly
- |
  woomera
- |
  woops
- |
  woozily
- |
  wooziness
- |
  woozy
- |
  Worcester
- |
  wordage
- |
  wordbook
- |
  wordily
- |
  wordiness
- |
  wording
- |
  wordless
- |
  wordlessly
- |
  wordplay
- |
  words
- |
  Wordsworth
- |
  wordy
- |
  workability
- |
  workable
- |
  workableness
- |
  workaday
- |
  workaholic
- |
  workbench
- |
  workbook
- |
  workday
- |
  worker
- |
  workfare
- |
  workforce
- |
  workhorse
- |
  workhouse
- |
  working
- |
  workingman
- |
  workings
- |
  workload
- |
  workman
- |
  workmanlike
- |
  workmanly
- |
  workmanship
- |
  workout
- |
  workplace
- |
  workroom
- |
  works
- |
  worksheet
- |
  workshop
- |
  workspace
- |
  workstation
- |
  worktable
- |
  workup
- |
  workweek
- |
  World
- |
  world
- |
  worldliness
- |
  worldling
- |
  worldly
- |
  worlds
- |
  worldview
- |
  worldwide
- |
  wormhole
- |
  worminess
- |
  worms
- |
  wormwood
- |
  wormy
- |
  worried
- |
  worriedly
- |
  worrier
- |
  worriment
- |
  worrisome
- |
  worry
- |
  worrying
- |
  worryingly
- |
  worrywart
- |
  worse
- |
  worsen
- |
  worsening
- |
  Worship
- |
  worship
- |
  worshiper
- |
  worshipful
- |
  worshipfully
- |
  worshipper
- |
  worst
- |
  worsted
- |
  worth
- |
  worthily
- |
  worthiness
- |
  worthless
- |
  worthwhile
- |
  worthy
- |
  would
- |
  wouldest
- |
  wouldst
- |
  wound
- |
  wounded
- |
  woven
- |
  wrack
- |
  wraith
- |
  wraithlike
- |
  Wrangell
- |
  wrangle
- |
  wrangler
- |
  wrangling
- |
  wraparound
- |
  wrapper
- |
  wrapping
- |
  wrappings
- |
  wrapt
- |
  wrasse
- |
  wrath
- |
  wrathful
- |
  wrathfully
- |
  wrathfulness
- |
  wreak
- |
  wreaker
- |
  wreath
- |
  wreathe
- |
  wreck
- |
  wreckage
- |
  wrecker
- |
  wrench
- |
  wrenching
- |
  wrest
- |
  wrester
- |
  wrestle
- |
  wrestler
- |
  wrestling
- |
  wretch
- |
  wretched
- |
  wretchedly
- |
  wretchedness
- |
  wrier
- |
  wriest
- |
  wriggle
- |
  wriggler
- |
  wriggly
- |
  Wright
- |
  wright
- |
  wring
- |
  wringer
- |
  wrinkle
- |
  wrinkled
- |
  wrinkly
- |
  wrist
- |
  wristband
- |
  wristlet
- |
  wristwatch
- |
  writable
- |
  write
- |
  writeable
- |
  writer
- |
  writhe
- |
  writing
- |
  Writings
- |
  writings
- |
  written
- |
  Wroclaw
- |
  wrong
- |
  wrongdoer
- |
  wrongdoing
- |
  wrongful
- |
  wrongfully
- |
  wrongfulness
- |
  wrongheaded
- |
  wrongly
- |
  wrongness
- |
  wrote
- |
  wroth
- |
  wrought
- |
  wrung
- |
  wryly
- |
  wryneck
- |
  wryness
- |
  Wuhan
- |
  wunderkind
- |
  wunderkinder
- |
  Wuppertal
- |
  wurst
- |
  Wusih
- |
  wussy
- |
  Wyandot
- |
  Wyandotte
- |
  Wyatt
- |
  Wycherley
- |
  Wycliffe
- |
  Wyeth
- |
  Wylie
- |
  Wyoming
- |
  Wyomingite
- |
  WYSIWYG
- |
  wysiwyg
- |
  Xanadu
- |
  Xanthippe
- |
  Xanthus
- |
  Xantippe
- |
  Xavier
- |
  xebec
- |
  xenon
- |
  Xenophanes
- |
  xenophobe
- |
  xenophobia
- |
  xenophobic
- |
  Xenophon
- |
  xeric
- |
  xerographic
- |
  xerography
- |
  xerophyte
- |
  xerophytic
- |
  Xerox
- |
  xerox
- |
  Xerxes
- |
  Xhosa
- |
  Xiamen
- |
  Xingu
- |
  Xizang
- |
  Xuzhou
- |
  xylem
- |
  xyloid
- |
  xylophone
- |
  xylophonist
- |
  yacht
- |
  yachting
- |
  yachtsman
- |
  yachtswoman
- |
  Yahoo
- |
  yahoo
- |
  Yahveh
- |
  Yahwe
- |
  Yahweh
- |
  Yakima
- |
  Yalta
- |
  yammer
- |
  yammerer
- |
  Yamoussoukro
- |
  Yamuna
- |
  Yangon
- |
  Yangtze
- |
  Yankee
- |
  yanqui
- |
  Yaounde
- |
  yapper
- |
  yappy
- |
  Yaqui
- |
  yardage
- |
  yardarm
- |
  yardman
- |
  yardmaster
- |
  yardstick
- |
  Yaren
- |
  yarmelke
- |
  yarmulka
- |
  yarmulke
- |
  Yaroslavl
- |
  yarrow
- |
  yawner
- |
  yawper
- |
  Yazoo
- |
  ycleped
- |
  yclept
- |
  yearbook
- |
  yearling
- |
  yearlong
- |
  yearly
- |
  yearn
- |
  yearning
- |
  years
- |
  yeast
- |
  yeasty
- |
  Yeats
- |
  Yeatsian
- |
  Yellow
- |
  yellow
- |
  yellowish
- |
  Yellowknife
- |
  yellowness
- |
  Yellowstone
- |
  yellowy
- |
  Yeltsin
- |
  Yemen
- |
  Yemeni
- |
  Yemenite
- |
  Yenisei
- |
  Yenisey
- |
  yenta
- |
  yeoman
- |
  yeomanly
- |
  yeomanry
- |
  Yerevan
- |
  yeshiva
- |
  yeshivah
- |
  yeshivoth
- |
  yester
- |
  yesterday
- |
  yesterdays
- |
  yesteryear
- |
  Yevtushenko
- |
  Yiddish
- |
  yield
- |
  yielding
- |
  yikes
- |
  yippee
- |
  yippie
- |
  yodel
- |
  yodeler
- |
  yodeller
- |
  yoghurt
- |
  yogic
- |
  yogin
- |
  yogurt
- |
  yokel
- |
  yokes
- |
  Yokohama
- |
  Yokosuka
- |
  Yolanda
- |
  yolked
- |
  yonder
- |
  Yonkers
- |
  Yorkie
- |
  Yorkshire
- |
  Yorktown
- |
  Yoruba
- |
  Yoruban
- |
  Yosemite
- |
  Young
- |
  young
- |
  youngish
- |
  youngling
- |
  youngster
- |
  Youngstown
- |
  yours
- |
  yourself
- |
  yourselves
- |
  youth
- |
  youthful
- |
  youthfully
- |
  youthfulness
- |
  ytterbium
- |
  yttrium
- |
  Yucatan
- |
  yucca
- |
  yucky
- |
  Yugoslav
- |
  Yugoslavia
- |
  Yugoslavian
- |
  Yukon
- |
  Yuletide
- |
  yuletide
- |
  yummy
- |
  Yupik
- |
  yuppie
- |
  yuppiedom
- |
  yuppify
- |
  yuppy
- |
  Yvette
- |
  Yvonne
- |
  Zacatecas
- |
  Zachariah
- |
  Zacharias
- |
  Zachary
- |
  zaftig
- |
  Zagreb
- |
  Zaharias
- |
  Zaire
- |
  zaire
- |
  Zairean
- |
  Zairian
- |
  Zambesi
- |
  Zambezi
- |
  Zambia
- |
  Zambian
- |
  zanily
- |
  zaniness
- |
  Zanzibar
- |
  Zapata
- |
  Zapopan
- |
  Zaporozhye
- |
  zapper
- |
  Zaragoza
- |
  Zarathustra
- |
  Zarqa
- |
  zazen
- |
  Zealot
- |
  zealot
- |
  zealotry
- |
  zealous
- |
  zealously
- |
  zealousness
- |
  zebra
- |
  Zechariah
- |
  Zedekiah
- |
  Zedong
- |
  Zeitgeist
- |
  zeitgeist
- |
  Zelda
- |
  zenana
- |
  Zenger
- |
  zenith
- |
  zenithal
- |
  zeolite
- |
  Zephaniah
- |
  Zephyr
- |
  zephyr
- |
  Zephyrus
- |
  Zeppelin
- |
  zeppelin
- |
  zestful
- |
  zestfully
- |
  zestfulness
- |
  zesty
- |
  Zetland
- |
  zeugma
- |
  zeugmatic
- |
  Zhangjiakou
- |
  Zhdanov
- |
  Zhengzhou
- |
  Zhukov
- |
  zidovudine
- |
  Ziegfeld
- |
  ziggurat
- |
  zigzag
- |
  zilch
- |
  zillion
- |
  Zimbabwe
- |
  Zimbabwean
- |
  zinfandel
- |
  zinger
- |
  zingy
- |
  zinnia
- |
  Zionism
- |
  Zionist
- |
  zipper
- |
  zippy
- |
  zircon
- |
  zirconium
- |
  zither
- |
  zitherist
- |
  zloty
- |
  zodiac
- |
  zodiacal
- |
  zoftig
- |
  Zomba
- |
  zombi
- |
  zombie
- |
  zombielike
- |
  zonal
- |
  zonally
- |
  zoned
- |
  zoning
- |
  zonked
- |
  zoogeography
- |
  zookeeper
- |
  zoologic
- |
  zoological
- |
  zoologist
- |
  zoology
- |
  zoomorphic
- |
  zoomorphism
- |
  zoophyte
- |
  zoophytic
- |
  zooplankton
- |
  zoospore
- |
  zootsuiter
- |
  Zoroaster
- |
  Zoroastrian
- |
  Zouave
- |
  zounds
- |
  zoysia
- |
  zucchetto
- |
  zucchini
- |
  Zululand
- |
  Zurich
- |
  zwieback
- |
  Zwingli
- |
  Zwinglian
- |
  zydeco
- |
  zygoses
- |
  zygosis
- |
  zygote
- |
  zygotic
- |
  zymurgy
word_to_guess:
- p
- a
- m
- p
- l
- o
- n
- a
